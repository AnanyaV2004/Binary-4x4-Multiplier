.INCLUDE TSMC_180nm.txt
* .include 22nm_MGK.pm
* .OPTIONS GMIN=1e-20 
* .option POST
* .options ABSTOL=1e-18 

.PARAM X=180n
.PARAM tr=10
.PARAM Src_Voltage = 1
.temp 25
.global GND 

*******Supply********
Vdd VDD GND dc= 'Src_Voltage'

**********SUBCKT AND*********
.SUBCKT and nodeA nodeB nodeOut node1 GND

* * ****Capacitive Load*********
* Cout nodeOut GND 0.001f
*M1 Drain Gate Source Body The name of model used in the model file included
Mp1 node5 nodeA node1 node1 pmos W={2*X} L={X}
Mp2 node5 nodeB node1 node1 pmos W={2*X} L={X}
Mn1 node4 nodeA GND GND nmos W={2*X} L={X}
Mn2 node5 nodeB node4 GND nmos W={2*X} L={X}
Mp3 nodeOut node5 node1 node1 pmos W={2*X} L={X}
Mn3 nodeOut node5 GND GND nmos W={2*X} L={X}

.ENDS and

**********SUBCKT INVERTER*********
.SUBCKT inv input output VDD GND

*M1 Drain Gate Source Body The name of model used in the model file included
Mp output input VDD VDD pmos W={2*X} L={X}
Mn output input GND GND nmos W={2*X} L={X}

.ENDS inv

**********SUBCKT XOR*********
.SUBCKT xor A B OUT VDD GND

XN1 A A_ VDD GND inv
XN2 B B_ VDD GND inv

*M1 Drain Gate Source Body The name of model used in the model file included
Mn1 node1 A_ GND GND nmos W={2*X} L={X}
Mn2 OUT B_ node1 GND nmos W={2*X} L={X}
Mn3 OUT B node2 GND nmos W={2*X} L={X}
Mn4 node2 A GND GND nmos W={2*X} L={X}

Mp1 OUT A_ node3 VDD pmos W={2*X} L={X}
Mp2 node3 B VDD VDD pmos W={2*X} L={X}
Mp3 node4 B_ VDD VDD pmos W={2*X} L={X}
Mp4 OUT A node4 VDD pmos W={2*X} L={X}

.ENDS xor

**********SUBCKT HALF ADDER*********
.SUBCKT halfadder A B VDD GND SUM CARRY

XH1 A B SUM VDD GND xor
XH2 A B CARRY VDD GND and

.ENDS halfadder


**********OR GATE*********
.SUBCKT or A B OUT VDD GND

*M1 Drain Gate Source Body The name of model used in the model file included
Mp1 node5 B TMP VDD pmos W={2*X} L={X}
Mp2 TMP A VDD VDD pmos W={2*X} L={X}
Mn1 node5 A GND GND nmos W={2*X} L={X}
Mn2 node5 B GND GND nmos W={2*X} L={X}
Mp3 OUT node5 VDD VDD pmos W={2*X} L={X}
Mn3 OUT node5 GND GND nmos W={2*X} L={X}

.ENDS or


**********SUBCKT FULL ADDER*********
.SUBCKT full_adder A B C SUM CARRY VDD GND
 XW1 A B VDD GND S0 C0 halfadder
 XW2 S0 C SUM VDD GND xor
 XW3 S0 C TMP VDD GND and
 XW4 C0 TMP CARRY VDD GND or
.ENDS full_adder


************** MAIN CIRCUIT MULTIPLIER ****************
*******************************************************

******AND GATES LEVELS********************
 XA1 A3 B3 O1 VDD GND and
 XA2 A3 B2 O2 VDD GND and
 XA3 A2 B3 O3 VDD GND and
 XA4 A1 B3 O4 VDD GND and
 XA5 A3 B1 O5 VDD GND and
 XA6 A2 B2 O6 VDD GND and
 XA7 A2 B1 O7 VDD GND and
 XA8 A3 B0 O8 VDD GND and
 XA9 A0 B3 O9 VDD GND and
 XA10 A1 B2 O10 VDD GND and
 XA11 A1 B1 O11 VDD GND and
 XA12 A2 B0 O12 VDD GND and
 XA13 A0 B2 O13 VDD GND and
 XA14 A1 B0 O14 VDD GND and
 XA15 A0 B1 O15 VDD GND and
 XA16 A0 B0 P0 VDD GND and
 *****************************************


 *************NEXT ADDER PART*************
* full_adder A B C SUM CARRY VDD GND
* halfadder A B VDD GND SUM CARRY

 XFA1 O2 O3 M1 L2 L1 VDD GND full_adder
 XHA2 O7 O8 VDD GND L4 L3 halfadder
 XHA3 O11 O12 VDD GND L6 L5 halfadder
 XHA4 O14 O15 VDD GND P1 L7 halfadder
 XFA5 O1 L1 M7 P6 C5 VDD GND full_adder
 XFA6 O5 O6 L3 M2 M1 VDD GND full_adder
 XFA7 L4 O10 L5 M4 M3 VDD GND full_adder
 XFA8 L6 O13 L7 P2 M5 VDD GND full_adder 
 XFA9 L2 M8 M10 P5 M7 VDD GND full_adder
 XFA10 O4 M2 M3 M9 M8 VDD GND full_adder
 XHA11 M9 M11 VDD GND P4 M10 halfadder
 XFA12 O9 M4 M5 P3 M11 VDD GND full_adder

******************************************


*********PROPAGATION DELAYS*********

VinA0 A3 GND PWL (0 0 {100} 0 {100+tr} 1)
VinA1 A2 GND PWL (0 0 {100} 0 {100+tr} 0)
VinA2 A1 GND PWL (0 0 {100} 0 {100+tr} 1)
VinA3 A0 GND PWL (0 0 {100} 0 {100+tr} 1)
VinB0 B3 GND PWL (0 0 {100} 0 {100+tr} 1)
VinB1 B2 GND PWL (0 0 {100} 0 {100+tr} 0)
VinB2 B1 GND PWL (0 0 {100} 0 {100+tr} 1)
VinB3 B0 GND PWL (0 0 {100} 0 {100+tr} 0)

***********DELAY*****************
.tran 0.1 100000

.control
run 
meas tran delay trig v(A0) val=0.5 rise=1 targ v(P6) val=0.5 rise=1

echo "(1,0,1,1,1,0,1,0)             $&delay" >> delay.txt
.endc 

.end


