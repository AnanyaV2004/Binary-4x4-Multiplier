magic
tech scmos
timestamp 1669632834
<< nwell >>
rect 45 -823 68 -748
rect 105 -823 128 -748
rect 165 -823 188 -748
rect 225 -823 248 -748
rect 285 -823 308 -748
rect 345 -823 368 -748
rect 405 -823 428 -748
rect 465 -823 488 -748
rect 525 -823 548 -748
rect 585 -823 608 -748
rect 645 -823 668 -748
rect 705 -823 728 -748
rect 765 -823 788 -748
rect 825 -823 848 -748
rect 885 -823 908 -748
rect 945 -823 968 -748
rect 22 -963 45 -888
rect 132 -906 155 -881
rect 132 -1042 155 -917
rect 367 -943 390 -868
rect 477 -886 500 -861
rect 477 -1022 500 -897
rect 604 -947 627 -872
rect 714 -890 737 -865
rect 714 -1026 737 -901
rect 787 -947 810 -872
rect 897 -890 920 -865
rect 897 -1026 920 -901
rect 65 -1154 88 -1079
rect 166 -1097 189 -1072
rect 53 -1248 76 -1174
rect 166 -1233 189 -1108
rect -242 -1513 -219 -1438
rect -132 -1456 -109 -1431
rect -132 -1592 -109 -1467
rect 187 -1512 210 -1437
rect 297 -1455 320 -1430
rect 297 -1591 320 -1466
rect 416 -1512 439 -1437
rect 526 -1455 549 -1430
rect 526 -1591 549 -1466
rect 655 -1509 678 -1434
rect 765 -1452 788 -1427
rect 765 -1588 788 -1463
rect -199 -1704 -176 -1629
rect -98 -1647 -75 -1622
rect -211 -1799 -188 -1724
rect -98 -1783 -75 -1658
rect 230 -1703 253 -1628
rect 331 -1646 354 -1621
rect 218 -1798 241 -1723
rect 331 -1782 354 -1657
rect 459 -1703 482 -1628
rect 560 -1646 583 -1621
rect 447 -1798 470 -1723
rect 560 -1782 583 -1657
rect 698 -1700 721 -1625
rect 799 -1643 822 -1618
rect 686 -1795 709 -1720
rect 799 -1779 822 -1654
rect -45 -1991 -22 -1916
rect 65 -1934 88 -1909
rect 65 -2070 88 -1945
rect 193 -1991 216 -1916
rect 303 -1934 326 -1909
rect 303 -2070 326 -1945
rect 437 -1980 460 -1905
rect 547 -1923 570 -1898
rect 547 -2059 570 -1934
rect 630 -1988 653 -1913
rect 740 -1931 763 -1906
rect 740 -2067 763 -1942
rect -2 -2182 21 -2107
rect 99 -2125 122 -2100
rect -14 -2277 9 -2202
rect 99 -2261 122 -2136
rect 236 -2182 259 -2107
rect 337 -2125 360 -2100
rect 224 -2277 247 -2202
rect 337 -2261 360 -2136
rect 673 -2179 696 -2104
rect 774 -2122 797 -2097
rect 661 -2274 684 -2199
rect 774 -2258 797 -2133
<< ntransistor >>
rect 20 -761 24 -759
rect 80 -761 84 -759
rect 140 -761 144 -759
rect 200 -761 204 -759
rect 260 -761 264 -759
rect 320 -761 324 -759
rect 380 -761 384 -759
rect 440 -761 444 -759
rect 500 -761 504 -759
rect 560 -761 564 -759
rect 620 -761 624 -759
rect 680 -761 684 -759
rect 740 -761 744 -759
rect 800 -761 804 -759
rect 860 -761 864 -759
rect 920 -761 924 -759
rect 20 -786 24 -784
rect 80 -786 84 -784
rect 140 -786 144 -784
rect 200 -786 204 -784
rect 260 -786 264 -784
rect 320 -786 324 -784
rect 380 -786 384 -784
rect 440 -786 444 -784
rect 500 -786 504 -784
rect 560 -786 564 -784
rect 620 -786 624 -784
rect 680 -786 684 -784
rect 740 -786 744 -784
rect 800 -786 804 -784
rect 860 -786 864 -784
rect 920 -786 924 -784
rect 20 -811 24 -809
rect 80 -811 84 -809
rect 140 -811 144 -809
rect 200 -811 204 -809
rect 260 -811 264 -809
rect 320 -811 324 -809
rect 380 -811 384 -809
rect 440 -811 444 -809
rect 500 -811 504 -809
rect 560 -811 564 -809
rect 620 -811 624 -809
rect 680 -811 684 -809
rect 740 -811 744 -809
rect 800 -811 804 -809
rect 860 -811 864 -809
rect 920 -811 924 -809
rect 416 -874 420 -872
rect 653 -878 657 -876
rect 836 -878 840 -876
rect 342 -881 346 -879
rect 579 -885 583 -883
rect 762 -885 766 -883
rect 71 -894 75 -892
rect -3 -901 1 -899
rect 342 -906 346 -904
rect 452 -910 456 -908
rect 579 -910 583 -908
rect 762 -910 766 -908
rect 689 -914 693 -912
rect 872 -914 876 -912
rect -3 -926 1 -924
rect 107 -930 111 -928
rect 342 -931 346 -929
rect 416 -935 420 -933
rect 579 -935 583 -933
rect 762 -935 766 -933
rect 653 -939 657 -937
rect 836 -939 840 -937
rect -3 -951 1 -949
rect 71 -955 75 -953
rect 416 -960 420 -958
rect 653 -964 657 -962
rect 836 -964 840 -962
rect 71 -980 75 -978
rect 452 -985 456 -983
rect 689 -989 693 -987
rect 872 -989 876 -987
rect 107 -1005 111 -1003
rect 416 -1010 420 -1008
rect 653 -1014 657 -1012
rect 836 -1014 840 -1012
rect 71 -1030 75 -1028
rect 105 -1085 109 -1083
rect 40 -1092 44 -1090
rect 40 -1117 44 -1115
rect 141 -1121 145 -1119
rect 40 -1142 44 -1140
rect 105 -1146 109 -1144
rect 105 -1171 109 -1169
rect 15 -1187 19 -1185
rect 141 -1196 145 -1194
rect 15 -1212 19 -1210
rect 105 -1221 109 -1219
rect 28 -1237 32 -1235
rect 704 -1440 708 -1438
rect -193 -1444 -189 -1442
rect 236 -1443 240 -1441
rect 465 -1443 469 -1441
rect 630 -1447 634 -1445
rect -267 -1451 -263 -1449
rect 162 -1450 166 -1448
rect 391 -1450 395 -1448
rect -267 -1476 -263 -1474
rect 162 -1475 166 -1473
rect -157 -1480 -153 -1478
rect 630 -1472 634 -1470
rect 391 -1475 395 -1473
rect 272 -1479 276 -1477
rect 740 -1476 744 -1474
rect 501 -1479 505 -1477
rect -267 -1501 -263 -1499
rect 162 -1500 166 -1498
rect -193 -1505 -189 -1503
rect 630 -1497 634 -1495
rect 391 -1500 395 -1498
rect 236 -1504 240 -1502
rect 704 -1501 708 -1499
rect 465 -1504 469 -1502
rect 704 -1526 708 -1524
rect -193 -1530 -189 -1528
rect 236 -1529 240 -1527
rect 465 -1529 469 -1527
rect 740 -1551 744 -1549
rect -157 -1555 -153 -1553
rect 272 -1554 276 -1552
rect 501 -1554 505 -1552
rect 704 -1576 708 -1574
rect -193 -1580 -189 -1578
rect 236 -1579 240 -1577
rect 465 -1579 469 -1577
rect 738 -1631 742 -1629
rect -159 -1635 -155 -1633
rect 270 -1634 274 -1632
rect 499 -1634 503 -1632
rect 673 -1638 677 -1636
rect -224 -1642 -220 -1640
rect 205 -1641 209 -1639
rect 434 -1641 438 -1639
rect -224 -1667 -220 -1665
rect 205 -1666 209 -1664
rect -123 -1671 -119 -1669
rect 673 -1663 677 -1661
rect 434 -1666 438 -1664
rect 306 -1670 310 -1668
rect 774 -1667 778 -1665
rect 535 -1670 539 -1668
rect -224 -1692 -220 -1690
rect 205 -1691 209 -1689
rect -159 -1696 -155 -1694
rect 673 -1688 677 -1686
rect 434 -1691 438 -1689
rect 270 -1695 274 -1693
rect 738 -1692 742 -1690
rect 499 -1695 503 -1693
rect 738 -1717 742 -1715
rect -159 -1721 -155 -1719
rect 270 -1720 274 -1718
rect 499 -1720 503 -1718
rect 648 -1733 652 -1731
rect -249 -1737 -245 -1735
rect 180 -1736 184 -1734
rect 409 -1736 413 -1734
rect 774 -1742 778 -1740
rect -123 -1746 -119 -1744
rect 306 -1745 310 -1743
rect 535 -1745 539 -1743
rect 648 -1758 652 -1756
rect -249 -1762 -245 -1760
rect 180 -1761 184 -1759
rect 409 -1761 413 -1759
rect 738 -1767 742 -1765
rect -159 -1771 -155 -1769
rect 270 -1770 274 -1768
rect 499 -1770 503 -1768
rect 661 -1783 665 -1781
rect -236 -1787 -232 -1785
rect 193 -1786 197 -1784
rect 422 -1786 426 -1784
rect 486 -1911 490 -1909
rect 412 -1918 416 -1916
rect 4 -1922 8 -1920
rect 242 -1922 246 -1920
rect 679 -1919 683 -1917
rect 605 -1926 609 -1924
rect -70 -1929 -66 -1927
rect 168 -1929 172 -1927
rect 412 -1943 416 -1941
rect -70 -1954 -66 -1952
rect 522 -1947 526 -1945
rect 168 -1954 172 -1952
rect 40 -1958 44 -1956
rect 605 -1951 609 -1949
rect 715 -1955 719 -1953
rect 278 -1958 282 -1956
rect 412 -1968 416 -1966
rect -70 -1979 -66 -1977
rect 486 -1972 490 -1970
rect 168 -1979 172 -1977
rect 4 -1983 8 -1981
rect 605 -1976 609 -1974
rect 679 -1980 683 -1978
rect 242 -1983 246 -1981
rect 486 -1997 490 -1995
rect 679 -2005 683 -2003
rect 4 -2008 8 -2006
rect 242 -2008 246 -2006
rect 522 -2022 526 -2020
rect 715 -2030 719 -2028
rect 40 -2033 44 -2031
rect 278 -2033 282 -2031
rect 486 -2047 490 -2045
rect 679 -2055 683 -2053
rect 4 -2058 8 -2056
rect 242 -2058 246 -2056
rect 713 -2110 717 -2108
rect 38 -2113 42 -2111
rect 276 -2113 280 -2111
rect 648 -2117 652 -2115
rect -27 -2120 -23 -2118
rect 211 -2120 215 -2118
rect -27 -2145 -23 -2143
rect 648 -2142 652 -2140
rect 211 -2145 215 -2143
rect 74 -2149 78 -2147
rect 749 -2146 753 -2144
rect 312 -2149 316 -2147
rect -27 -2170 -23 -2168
rect 648 -2167 652 -2165
rect 211 -2170 215 -2168
rect 38 -2174 42 -2172
rect 713 -2171 717 -2169
rect 276 -2174 280 -2172
rect 713 -2196 717 -2194
rect 38 -2199 42 -2197
rect 276 -2199 280 -2197
rect 623 -2212 627 -2210
rect -52 -2215 -48 -2213
rect 186 -2215 190 -2213
rect 749 -2221 753 -2219
rect 74 -2224 78 -2222
rect 312 -2224 316 -2222
rect 623 -2237 627 -2235
rect -52 -2240 -48 -2238
rect 186 -2240 190 -2238
rect 713 -2246 717 -2244
rect 38 -2249 42 -2247
rect 276 -2249 280 -2247
rect 636 -2262 640 -2260
rect -39 -2265 -35 -2263
rect 199 -2265 203 -2263
<< ptransistor >>
rect 51 -761 59 -759
rect 111 -761 119 -759
rect 171 -761 179 -759
rect 231 -761 239 -759
rect 291 -761 299 -759
rect 351 -761 359 -759
rect 411 -761 419 -759
rect 471 -761 479 -759
rect 531 -761 539 -759
rect 591 -761 599 -759
rect 651 -761 659 -759
rect 711 -761 719 -759
rect 771 -761 779 -759
rect 831 -761 839 -759
rect 891 -761 899 -759
rect 951 -761 959 -759
rect 51 -786 59 -784
rect 111 -786 119 -784
rect 171 -786 179 -784
rect 231 -786 239 -784
rect 291 -786 299 -784
rect 351 -786 359 -784
rect 411 -786 419 -784
rect 471 -786 479 -784
rect 531 -786 539 -784
rect 591 -786 599 -784
rect 651 -786 659 -784
rect 711 -786 719 -784
rect 771 -786 779 -784
rect 831 -786 839 -784
rect 891 -786 899 -784
rect 951 -786 959 -784
rect 51 -811 59 -809
rect 111 -811 119 -809
rect 171 -811 179 -809
rect 231 -811 239 -809
rect 291 -811 299 -809
rect 351 -811 359 -809
rect 411 -811 419 -809
rect 471 -811 479 -809
rect 531 -811 539 -809
rect 591 -811 599 -809
rect 651 -811 659 -809
rect 711 -811 719 -809
rect 771 -811 779 -809
rect 831 -811 839 -809
rect 891 -811 899 -809
rect 951 -811 959 -809
rect 483 -874 491 -872
rect 720 -878 728 -876
rect 903 -878 911 -876
rect 373 -881 381 -879
rect 610 -885 618 -883
rect 793 -885 801 -883
rect 138 -894 146 -892
rect 28 -901 36 -899
rect 373 -906 381 -904
rect 483 -910 491 -908
rect 610 -910 618 -908
rect 793 -910 801 -908
rect 720 -914 728 -912
rect 903 -914 911 -912
rect 28 -926 36 -924
rect 138 -930 146 -928
rect 373 -931 381 -929
rect 483 -935 491 -933
rect 610 -935 618 -933
rect 793 -935 801 -933
rect 720 -939 728 -937
rect 903 -939 911 -937
rect 28 -951 36 -949
rect 138 -955 146 -953
rect 483 -960 491 -958
rect 720 -964 728 -962
rect 903 -964 911 -962
rect 138 -980 146 -978
rect 483 -985 491 -983
rect 720 -989 728 -987
rect 903 -989 911 -987
rect 138 -1005 146 -1003
rect 483 -1010 491 -1008
rect 720 -1014 728 -1012
rect 903 -1014 911 -1012
rect 138 -1030 146 -1028
rect 172 -1085 180 -1083
rect 71 -1092 79 -1090
rect 71 -1117 79 -1115
rect 172 -1121 180 -1119
rect 71 -1142 79 -1140
rect 172 -1146 180 -1144
rect 172 -1171 180 -1169
rect 59 -1187 67 -1185
rect 172 -1196 180 -1194
rect 59 -1212 67 -1210
rect 172 -1221 180 -1219
rect 59 -1237 67 -1235
rect 771 -1440 779 -1438
rect -126 -1444 -118 -1442
rect 303 -1443 311 -1441
rect 532 -1443 540 -1441
rect 661 -1447 669 -1445
rect -236 -1451 -228 -1449
rect 193 -1450 201 -1448
rect 422 -1450 430 -1448
rect -236 -1476 -228 -1474
rect 193 -1475 201 -1473
rect -126 -1480 -118 -1478
rect 661 -1472 669 -1470
rect 422 -1475 430 -1473
rect 303 -1479 311 -1477
rect 771 -1476 779 -1474
rect 532 -1479 540 -1477
rect -236 -1501 -228 -1499
rect 193 -1500 201 -1498
rect -126 -1505 -118 -1503
rect 661 -1497 669 -1495
rect 422 -1500 430 -1498
rect 303 -1504 311 -1502
rect 771 -1501 779 -1499
rect 532 -1504 540 -1502
rect 771 -1526 779 -1524
rect -126 -1530 -118 -1528
rect 303 -1529 311 -1527
rect 532 -1529 540 -1527
rect 771 -1551 779 -1549
rect -126 -1555 -118 -1553
rect 303 -1554 311 -1552
rect 532 -1554 540 -1552
rect 771 -1576 779 -1574
rect -126 -1580 -118 -1578
rect 303 -1579 311 -1577
rect 532 -1579 540 -1577
rect 805 -1631 813 -1629
rect -92 -1635 -84 -1633
rect 337 -1634 345 -1632
rect 566 -1634 574 -1632
rect 704 -1638 712 -1636
rect -193 -1642 -185 -1640
rect 236 -1641 244 -1639
rect 465 -1641 473 -1639
rect -193 -1667 -185 -1665
rect 236 -1666 244 -1664
rect -92 -1671 -84 -1669
rect 704 -1663 712 -1661
rect 465 -1666 473 -1664
rect 337 -1670 345 -1668
rect 805 -1667 813 -1665
rect 566 -1670 574 -1668
rect -193 -1692 -185 -1690
rect 236 -1691 244 -1689
rect -92 -1696 -84 -1694
rect 704 -1688 712 -1686
rect 465 -1691 473 -1689
rect 337 -1695 345 -1693
rect 805 -1692 813 -1690
rect 566 -1695 574 -1693
rect 805 -1717 813 -1715
rect -92 -1721 -84 -1719
rect 337 -1720 345 -1718
rect 566 -1720 574 -1718
rect 692 -1733 700 -1731
rect -205 -1737 -197 -1735
rect 224 -1736 232 -1734
rect 453 -1736 461 -1734
rect 805 -1742 813 -1740
rect -92 -1746 -84 -1744
rect 337 -1745 345 -1743
rect 566 -1745 574 -1743
rect 692 -1758 700 -1756
rect -205 -1762 -197 -1760
rect 224 -1761 232 -1759
rect 453 -1761 461 -1759
rect 805 -1767 813 -1765
rect -92 -1771 -84 -1769
rect 337 -1770 345 -1768
rect 566 -1770 574 -1768
rect 692 -1783 700 -1781
rect -205 -1787 -197 -1785
rect 224 -1786 232 -1784
rect 453 -1786 461 -1784
rect 553 -1911 561 -1909
rect 443 -1918 451 -1916
rect 71 -1922 79 -1920
rect 309 -1922 317 -1920
rect 746 -1919 754 -1917
rect 636 -1926 644 -1924
rect -39 -1929 -31 -1927
rect 199 -1929 207 -1927
rect 443 -1943 451 -1941
rect -39 -1954 -31 -1952
rect 553 -1947 561 -1945
rect 199 -1954 207 -1952
rect 71 -1958 79 -1956
rect 636 -1951 644 -1949
rect 746 -1955 754 -1953
rect 309 -1958 317 -1956
rect 443 -1968 451 -1966
rect -39 -1979 -31 -1977
rect 553 -1972 561 -1970
rect 199 -1979 207 -1977
rect 71 -1983 79 -1981
rect 636 -1976 644 -1974
rect 746 -1980 754 -1978
rect 309 -1983 317 -1981
rect 553 -1997 561 -1995
rect 746 -2005 754 -2003
rect 71 -2008 79 -2006
rect 309 -2008 317 -2006
rect 553 -2022 561 -2020
rect 746 -2030 754 -2028
rect 71 -2033 79 -2031
rect 309 -2033 317 -2031
rect 553 -2047 561 -2045
rect 746 -2055 754 -2053
rect 71 -2058 79 -2056
rect 309 -2058 317 -2056
rect 780 -2110 788 -2108
rect 105 -2113 113 -2111
rect 343 -2113 351 -2111
rect 679 -2117 687 -2115
rect 4 -2120 12 -2118
rect 242 -2120 250 -2118
rect 4 -2145 12 -2143
rect 679 -2142 687 -2140
rect 242 -2145 250 -2143
rect 105 -2149 113 -2147
rect 780 -2146 788 -2144
rect 343 -2149 351 -2147
rect 4 -2170 12 -2168
rect 679 -2167 687 -2165
rect 242 -2170 250 -2168
rect 105 -2174 113 -2172
rect 780 -2171 788 -2169
rect 343 -2174 351 -2172
rect 780 -2196 788 -2194
rect 105 -2199 113 -2197
rect 343 -2199 351 -2197
rect 667 -2212 675 -2210
rect -8 -2215 0 -2213
rect 230 -2215 238 -2213
rect 780 -2221 788 -2219
rect 105 -2224 113 -2222
rect 343 -2224 351 -2222
rect 667 -2237 675 -2235
rect -8 -2240 0 -2238
rect 230 -2240 238 -2238
rect 780 -2246 788 -2244
rect 105 -2249 113 -2247
rect 343 -2249 351 -2247
rect 667 -2262 675 -2260
rect -8 -2265 0 -2263
rect 230 -2265 238 -2263
<< ndiffusion >>
rect 20 -759 24 -758
rect 80 -759 84 -758
rect 140 -759 144 -758
rect 200 -759 204 -758
rect 260 -759 264 -758
rect 320 -759 324 -758
rect 380 -759 384 -758
rect 440 -759 444 -758
rect 500 -759 504 -758
rect 560 -759 564 -758
rect 620 -759 624 -758
rect 680 -759 684 -758
rect 740 -759 744 -758
rect 800 -759 804 -758
rect 860 -759 864 -758
rect 920 -759 924 -758
rect 20 -762 24 -761
rect 80 -762 84 -761
rect 140 -762 144 -761
rect 200 -762 204 -761
rect 260 -762 264 -761
rect 320 -762 324 -761
rect 380 -762 384 -761
rect 440 -762 444 -761
rect 500 -762 504 -761
rect 560 -762 564 -761
rect 620 -762 624 -761
rect 680 -762 684 -761
rect 740 -762 744 -761
rect 800 -762 804 -761
rect 860 -762 864 -761
rect 920 -762 924 -761
rect 20 -784 24 -783
rect 80 -784 84 -783
rect 140 -784 144 -783
rect 200 -784 204 -783
rect 260 -784 264 -783
rect 320 -784 324 -783
rect 380 -784 384 -783
rect 440 -784 444 -783
rect 500 -784 504 -783
rect 560 -784 564 -783
rect 620 -784 624 -783
rect 680 -784 684 -783
rect 740 -784 744 -783
rect 800 -784 804 -783
rect 860 -784 864 -783
rect 920 -784 924 -783
rect 20 -787 24 -786
rect 80 -787 84 -786
rect 140 -787 144 -786
rect 200 -787 204 -786
rect 260 -787 264 -786
rect 320 -787 324 -786
rect 380 -787 384 -786
rect 440 -787 444 -786
rect 500 -787 504 -786
rect 560 -787 564 -786
rect 620 -787 624 -786
rect 680 -787 684 -786
rect 740 -787 744 -786
rect 800 -787 804 -786
rect 860 -787 864 -786
rect 920 -787 924 -786
rect 20 -809 24 -808
rect 80 -809 84 -808
rect 140 -809 144 -808
rect 200 -809 204 -808
rect 260 -809 264 -808
rect 320 -809 324 -808
rect 380 -809 384 -808
rect 440 -809 444 -808
rect 500 -809 504 -808
rect 560 -809 564 -808
rect 620 -809 624 -808
rect 680 -809 684 -808
rect 740 -809 744 -808
rect 800 -809 804 -808
rect 860 -809 864 -808
rect 920 -809 924 -808
rect 20 -812 24 -811
rect 80 -812 84 -811
rect 140 -812 144 -811
rect 200 -812 204 -811
rect 260 -812 264 -811
rect 320 -812 324 -811
rect 380 -812 384 -811
rect 440 -812 444 -811
rect 500 -812 504 -811
rect 560 -812 564 -811
rect 620 -812 624 -811
rect 680 -812 684 -811
rect 740 -812 744 -811
rect 800 -812 804 -811
rect 860 -812 864 -811
rect 920 -812 924 -811
rect 416 -872 420 -871
rect 342 -879 346 -878
rect 416 -875 420 -874
rect 653 -876 657 -875
rect 836 -876 840 -875
rect 342 -882 346 -881
rect 579 -883 583 -882
rect 653 -879 657 -878
rect 762 -883 766 -882
rect 836 -879 840 -878
rect 579 -886 583 -885
rect 71 -892 75 -891
rect 762 -886 766 -885
rect -3 -899 1 -898
rect 71 -895 75 -894
rect -3 -902 1 -901
rect 342 -904 346 -903
rect 342 -907 346 -906
rect 452 -908 456 -907
rect 579 -908 583 -907
rect 452 -911 456 -910
rect 579 -911 583 -910
rect 689 -912 693 -911
rect 762 -908 766 -907
rect 762 -911 766 -910
rect 689 -915 693 -914
rect 872 -912 876 -911
rect 872 -915 876 -914
rect -3 -924 1 -923
rect -3 -927 1 -926
rect 107 -928 111 -927
rect 342 -929 346 -928
rect 107 -931 111 -930
rect 342 -932 346 -931
rect 416 -933 420 -932
rect 579 -933 583 -932
rect 416 -936 420 -935
rect 579 -936 583 -935
rect 653 -937 657 -936
rect 762 -933 766 -932
rect 762 -936 766 -935
rect 653 -940 657 -939
rect 836 -937 840 -936
rect 836 -940 840 -939
rect -3 -949 1 -948
rect -3 -952 1 -951
rect 71 -953 75 -952
rect 71 -956 75 -955
rect 416 -958 420 -957
rect 416 -961 420 -960
rect 653 -962 657 -961
rect 836 -962 840 -961
rect 653 -965 657 -964
rect 836 -965 840 -964
rect 71 -978 75 -977
rect 71 -981 75 -980
rect 452 -983 456 -982
rect 452 -986 456 -985
rect 689 -987 693 -986
rect 872 -987 876 -986
rect 689 -990 693 -989
rect 872 -990 876 -989
rect 107 -1003 111 -1002
rect 107 -1006 111 -1005
rect 416 -1008 420 -1007
rect 416 -1011 420 -1010
rect 653 -1012 657 -1011
rect 836 -1012 840 -1011
rect 653 -1015 657 -1014
rect 836 -1015 840 -1014
rect 71 -1028 75 -1027
rect 71 -1031 75 -1030
rect 105 -1083 109 -1082
rect 40 -1090 44 -1089
rect 105 -1086 109 -1085
rect 40 -1093 44 -1092
rect 40 -1115 44 -1114
rect 40 -1118 44 -1117
rect 141 -1119 145 -1118
rect 141 -1122 145 -1121
rect 40 -1140 44 -1139
rect 40 -1143 44 -1142
rect 105 -1144 109 -1143
rect 105 -1147 109 -1146
rect 105 -1169 109 -1168
rect 105 -1172 109 -1171
rect 15 -1185 19 -1184
rect 15 -1188 19 -1187
rect 141 -1194 145 -1193
rect 141 -1197 145 -1196
rect 15 -1210 19 -1209
rect 15 -1213 19 -1212
rect 105 -1219 109 -1218
rect 105 -1222 109 -1221
rect 28 -1235 32 -1234
rect 28 -1238 32 -1237
rect -193 -1442 -189 -1441
rect 236 -1441 240 -1440
rect 465 -1441 469 -1440
rect 704 -1438 708 -1437
rect -267 -1449 -263 -1448
rect -193 -1445 -189 -1444
rect 162 -1448 166 -1447
rect 236 -1444 240 -1443
rect 391 -1448 395 -1447
rect 465 -1444 469 -1443
rect 630 -1445 634 -1444
rect 704 -1441 708 -1440
rect 630 -1448 634 -1447
rect 162 -1451 166 -1450
rect -267 -1452 -263 -1451
rect 391 -1451 395 -1450
rect -267 -1474 -263 -1473
rect 162 -1473 166 -1472
rect -267 -1477 -263 -1476
rect -157 -1478 -153 -1477
rect 162 -1476 166 -1475
rect 272 -1477 276 -1476
rect 391 -1473 395 -1472
rect 630 -1470 634 -1469
rect 391 -1476 395 -1475
rect 272 -1480 276 -1479
rect -157 -1481 -153 -1480
rect 501 -1477 505 -1476
rect 630 -1473 634 -1472
rect 740 -1474 744 -1473
rect 740 -1477 744 -1476
rect 501 -1480 505 -1479
rect -267 -1499 -263 -1498
rect 162 -1498 166 -1497
rect -267 -1502 -263 -1501
rect -193 -1503 -189 -1502
rect 162 -1501 166 -1500
rect 236 -1502 240 -1501
rect 391 -1498 395 -1497
rect 630 -1495 634 -1494
rect 391 -1501 395 -1500
rect 236 -1505 240 -1504
rect -193 -1506 -189 -1505
rect 465 -1502 469 -1501
rect 630 -1498 634 -1497
rect 704 -1499 708 -1498
rect 704 -1502 708 -1501
rect 465 -1505 469 -1504
rect -193 -1528 -189 -1527
rect 236 -1527 240 -1526
rect 465 -1527 469 -1526
rect 704 -1524 708 -1523
rect 704 -1527 708 -1526
rect 236 -1530 240 -1529
rect -193 -1531 -189 -1530
rect 465 -1530 469 -1529
rect -157 -1553 -153 -1552
rect 272 -1552 276 -1551
rect 501 -1552 505 -1551
rect 740 -1549 744 -1548
rect 740 -1552 744 -1551
rect 272 -1555 276 -1554
rect -157 -1556 -153 -1555
rect 501 -1555 505 -1554
rect -193 -1578 -189 -1577
rect 236 -1577 240 -1576
rect 465 -1577 469 -1576
rect 704 -1574 708 -1573
rect 704 -1577 708 -1576
rect 236 -1580 240 -1579
rect -193 -1581 -189 -1580
rect 465 -1580 469 -1579
rect -159 -1633 -155 -1632
rect 270 -1632 274 -1631
rect 499 -1632 503 -1631
rect 738 -1629 742 -1628
rect -224 -1640 -220 -1639
rect -159 -1636 -155 -1635
rect 205 -1639 209 -1638
rect 270 -1635 274 -1634
rect 434 -1639 438 -1638
rect 499 -1635 503 -1634
rect 673 -1636 677 -1635
rect 738 -1632 742 -1631
rect 673 -1639 677 -1638
rect 205 -1642 209 -1641
rect -224 -1643 -220 -1642
rect 434 -1642 438 -1641
rect -224 -1665 -220 -1664
rect 205 -1664 209 -1663
rect -224 -1668 -220 -1667
rect -123 -1669 -119 -1668
rect 205 -1667 209 -1666
rect 306 -1668 310 -1667
rect 434 -1664 438 -1663
rect 673 -1661 677 -1660
rect 434 -1667 438 -1666
rect 306 -1671 310 -1670
rect -123 -1672 -119 -1671
rect 535 -1668 539 -1667
rect 673 -1664 677 -1663
rect 774 -1665 778 -1664
rect 774 -1668 778 -1667
rect 535 -1671 539 -1670
rect -224 -1690 -220 -1689
rect 205 -1689 209 -1688
rect -224 -1693 -220 -1692
rect -159 -1694 -155 -1693
rect 205 -1692 209 -1691
rect 270 -1693 274 -1692
rect 434 -1689 438 -1688
rect 673 -1686 677 -1685
rect 434 -1692 438 -1691
rect 270 -1696 274 -1695
rect -159 -1697 -155 -1696
rect 499 -1693 503 -1692
rect 673 -1689 677 -1688
rect 738 -1690 742 -1689
rect 738 -1693 742 -1692
rect 499 -1696 503 -1695
rect -159 -1719 -155 -1718
rect 270 -1718 274 -1717
rect 499 -1718 503 -1717
rect 738 -1715 742 -1714
rect 738 -1718 742 -1717
rect 270 -1721 274 -1720
rect -159 -1722 -155 -1721
rect 499 -1721 503 -1720
rect -249 -1735 -245 -1734
rect 180 -1734 184 -1733
rect 409 -1734 413 -1733
rect 648 -1731 652 -1730
rect 648 -1734 652 -1733
rect 180 -1737 184 -1736
rect -249 -1738 -245 -1737
rect -123 -1744 -119 -1743
rect 409 -1737 413 -1736
rect 306 -1743 310 -1742
rect 535 -1743 539 -1742
rect 774 -1740 778 -1739
rect 774 -1743 778 -1742
rect 306 -1746 310 -1745
rect -123 -1747 -119 -1746
rect 535 -1746 539 -1745
rect -249 -1760 -245 -1759
rect 180 -1759 184 -1758
rect 409 -1759 413 -1758
rect 648 -1756 652 -1755
rect 648 -1759 652 -1758
rect 180 -1762 184 -1761
rect -249 -1763 -245 -1762
rect -159 -1769 -155 -1768
rect 409 -1762 413 -1761
rect 270 -1768 274 -1767
rect 499 -1768 503 -1767
rect 738 -1765 742 -1764
rect 738 -1768 742 -1767
rect 270 -1771 274 -1770
rect -159 -1772 -155 -1771
rect 499 -1771 503 -1770
rect -236 -1785 -232 -1784
rect 193 -1784 197 -1783
rect 422 -1784 426 -1783
rect 661 -1781 665 -1780
rect 661 -1784 665 -1783
rect 193 -1787 197 -1786
rect -236 -1788 -232 -1787
rect 422 -1787 426 -1786
rect 486 -1909 490 -1908
rect 4 -1920 8 -1919
rect 242 -1920 246 -1919
rect 412 -1916 416 -1915
rect 486 -1912 490 -1911
rect 679 -1917 683 -1916
rect 412 -1919 416 -1918
rect -70 -1927 -66 -1926
rect 4 -1923 8 -1922
rect 168 -1927 172 -1926
rect 242 -1923 246 -1922
rect 605 -1924 609 -1923
rect 679 -1920 683 -1919
rect 605 -1927 609 -1926
rect -70 -1930 -66 -1929
rect 168 -1930 172 -1929
rect 412 -1941 416 -1940
rect 412 -1944 416 -1943
rect -70 -1952 -66 -1951
rect -70 -1955 -66 -1954
rect 40 -1956 44 -1955
rect 168 -1952 172 -1951
rect 522 -1945 526 -1944
rect 522 -1948 526 -1947
rect 168 -1955 172 -1954
rect 40 -1959 44 -1958
rect 278 -1956 282 -1955
rect 605 -1949 609 -1948
rect 605 -1952 609 -1951
rect 715 -1953 719 -1952
rect 715 -1956 719 -1955
rect 278 -1959 282 -1958
rect 412 -1966 416 -1965
rect 412 -1969 416 -1968
rect -70 -1977 -66 -1976
rect -70 -1980 -66 -1979
rect 4 -1981 8 -1980
rect 168 -1977 172 -1976
rect 486 -1970 490 -1969
rect 486 -1973 490 -1972
rect 168 -1980 172 -1979
rect 4 -1984 8 -1983
rect 242 -1981 246 -1980
rect 605 -1974 609 -1973
rect 605 -1977 609 -1976
rect 679 -1978 683 -1977
rect 679 -1981 683 -1980
rect 242 -1984 246 -1983
rect 486 -1995 490 -1994
rect 486 -1998 490 -1997
rect 4 -2006 8 -2005
rect 242 -2006 246 -2005
rect 679 -2003 683 -2002
rect 679 -2006 683 -2005
rect 4 -2009 8 -2008
rect 242 -2009 246 -2008
rect 522 -2020 526 -2019
rect 522 -2023 526 -2022
rect 40 -2031 44 -2030
rect 278 -2031 282 -2030
rect 715 -2028 719 -2027
rect 715 -2031 719 -2030
rect 40 -2034 44 -2033
rect 278 -2034 282 -2033
rect 486 -2045 490 -2044
rect 486 -2048 490 -2047
rect 4 -2056 8 -2055
rect 242 -2056 246 -2055
rect 679 -2053 683 -2052
rect 679 -2056 683 -2055
rect 4 -2059 8 -2058
rect 242 -2059 246 -2058
rect 38 -2111 42 -2110
rect 276 -2111 280 -2110
rect 713 -2108 717 -2107
rect -27 -2118 -23 -2117
rect 38 -2114 42 -2113
rect 211 -2118 215 -2117
rect 276 -2114 280 -2113
rect 648 -2115 652 -2114
rect 713 -2111 717 -2110
rect 648 -2118 652 -2117
rect -27 -2121 -23 -2120
rect 211 -2121 215 -2120
rect -27 -2143 -23 -2142
rect -27 -2146 -23 -2145
rect 74 -2147 78 -2146
rect 211 -2143 215 -2142
rect 648 -2140 652 -2139
rect 211 -2146 215 -2145
rect 74 -2150 78 -2149
rect 312 -2147 316 -2146
rect 648 -2143 652 -2142
rect 749 -2144 753 -2143
rect 749 -2147 753 -2146
rect 312 -2150 316 -2149
rect -27 -2168 -23 -2167
rect -27 -2171 -23 -2170
rect 38 -2172 42 -2171
rect 211 -2168 215 -2167
rect 648 -2165 652 -2164
rect 211 -2171 215 -2170
rect 38 -2175 42 -2174
rect 276 -2172 280 -2171
rect 648 -2168 652 -2167
rect 713 -2169 717 -2168
rect 713 -2172 717 -2171
rect 276 -2175 280 -2174
rect 38 -2197 42 -2196
rect 276 -2197 280 -2196
rect 713 -2194 717 -2193
rect 713 -2197 717 -2196
rect 38 -2200 42 -2199
rect 276 -2200 280 -2199
rect -52 -2213 -48 -2212
rect 186 -2213 190 -2212
rect 623 -2210 627 -2209
rect 623 -2213 627 -2212
rect -52 -2216 -48 -2215
rect 186 -2216 190 -2215
rect 74 -2222 78 -2221
rect 312 -2222 316 -2221
rect 749 -2219 753 -2218
rect 749 -2222 753 -2221
rect 74 -2225 78 -2224
rect 312 -2225 316 -2224
rect -52 -2238 -48 -2237
rect 186 -2238 190 -2237
rect 623 -2235 627 -2234
rect 623 -2238 627 -2237
rect -52 -2241 -48 -2240
rect 186 -2241 190 -2240
rect 38 -2247 42 -2246
rect 276 -2247 280 -2246
rect 713 -2244 717 -2243
rect 713 -2247 717 -2246
rect 38 -2250 42 -2249
rect 276 -2250 280 -2249
rect -39 -2263 -35 -2262
rect 199 -2263 203 -2262
rect 636 -2260 640 -2259
rect 636 -2263 640 -2262
rect -39 -2266 -35 -2265
rect 199 -2266 203 -2265
<< pdiffusion >>
rect 51 -759 59 -758
rect 111 -759 119 -758
rect 171 -759 179 -758
rect 231 -759 239 -758
rect 291 -759 299 -758
rect 351 -759 359 -758
rect 411 -759 419 -758
rect 471 -759 479 -758
rect 531 -759 539 -758
rect 591 -759 599 -758
rect 651 -759 659 -758
rect 711 -759 719 -758
rect 771 -759 779 -758
rect 831 -759 839 -758
rect 891 -759 899 -758
rect 951 -759 959 -758
rect 51 -762 59 -761
rect 111 -762 119 -761
rect 171 -762 179 -761
rect 231 -762 239 -761
rect 291 -762 299 -761
rect 351 -762 359 -761
rect 411 -762 419 -761
rect 471 -762 479 -761
rect 531 -762 539 -761
rect 591 -762 599 -761
rect 651 -762 659 -761
rect 711 -762 719 -761
rect 771 -762 779 -761
rect 831 -762 839 -761
rect 891 -762 899 -761
rect 951 -762 959 -761
rect 51 -784 59 -783
rect 111 -784 119 -783
rect 171 -784 179 -783
rect 231 -784 239 -783
rect 291 -784 299 -783
rect 351 -784 359 -783
rect 411 -784 419 -783
rect 471 -784 479 -783
rect 531 -784 539 -783
rect 591 -784 599 -783
rect 651 -784 659 -783
rect 711 -784 719 -783
rect 771 -784 779 -783
rect 831 -784 839 -783
rect 891 -784 899 -783
rect 951 -784 959 -783
rect 51 -787 59 -786
rect 111 -787 119 -786
rect 171 -787 179 -786
rect 231 -787 239 -786
rect 291 -787 299 -786
rect 351 -787 359 -786
rect 411 -787 419 -786
rect 471 -787 479 -786
rect 531 -787 539 -786
rect 591 -787 599 -786
rect 651 -787 659 -786
rect 711 -787 719 -786
rect 771 -787 779 -786
rect 831 -787 839 -786
rect 891 -787 899 -786
rect 951 -787 959 -786
rect 51 -809 59 -808
rect 111 -809 119 -808
rect 171 -809 179 -808
rect 231 -809 239 -808
rect 291 -809 299 -808
rect 351 -809 359 -808
rect 411 -809 419 -808
rect 471 -809 479 -808
rect 531 -809 539 -808
rect 591 -809 599 -808
rect 651 -809 659 -808
rect 711 -809 719 -808
rect 771 -809 779 -808
rect 831 -809 839 -808
rect 891 -809 899 -808
rect 951 -809 959 -808
rect 51 -812 59 -811
rect 111 -812 119 -811
rect 171 -812 179 -811
rect 231 -812 239 -811
rect 291 -812 299 -811
rect 351 -812 359 -811
rect 411 -812 419 -811
rect 471 -812 479 -811
rect 531 -812 539 -811
rect 591 -812 599 -811
rect 651 -812 659 -811
rect 711 -812 719 -811
rect 771 -812 779 -811
rect 831 -812 839 -811
rect 891 -812 899 -811
rect 951 -812 959 -811
rect 483 -872 491 -871
rect 373 -879 381 -878
rect 483 -875 491 -874
rect 720 -876 728 -875
rect 903 -876 911 -875
rect 373 -882 381 -881
rect 610 -883 618 -882
rect 720 -879 728 -878
rect 793 -883 801 -882
rect 903 -879 911 -878
rect 610 -886 618 -885
rect 793 -886 801 -885
rect 138 -892 146 -891
rect 28 -899 36 -898
rect 138 -895 146 -894
rect 28 -902 36 -901
rect 373 -904 381 -903
rect 373 -907 381 -906
rect 483 -908 491 -907
rect 610 -908 618 -907
rect 483 -911 491 -910
rect 610 -911 618 -910
rect 793 -908 801 -907
rect 720 -912 728 -911
rect 720 -915 728 -914
rect 793 -911 801 -910
rect 903 -912 911 -911
rect 903 -915 911 -914
rect 28 -924 36 -923
rect 28 -927 36 -926
rect 138 -928 146 -927
rect 373 -929 381 -928
rect 138 -931 146 -930
rect 373 -932 381 -931
rect 483 -933 491 -932
rect 610 -933 618 -932
rect 483 -936 491 -935
rect 610 -936 618 -935
rect 793 -933 801 -932
rect 720 -937 728 -936
rect 720 -940 728 -939
rect 793 -936 801 -935
rect 903 -937 911 -936
rect 903 -940 911 -939
rect 28 -949 36 -948
rect 28 -952 36 -951
rect 138 -953 146 -952
rect 138 -956 146 -955
rect 483 -958 491 -957
rect 483 -961 491 -960
rect 720 -962 728 -961
rect 903 -962 911 -961
rect 720 -965 728 -964
rect 903 -965 911 -964
rect 138 -978 146 -977
rect 138 -981 146 -980
rect 483 -983 491 -982
rect 483 -986 491 -985
rect 720 -987 728 -986
rect 903 -987 911 -986
rect 720 -990 728 -989
rect 903 -990 911 -989
rect 138 -1003 146 -1002
rect 138 -1006 146 -1005
rect 483 -1008 491 -1007
rect 483 -1011 491 -1010
rect 720 -1012 728 -1011
rect 903 -1012 911 -1011
rect 720 -1015 728 -1014
rect 903 -1015 911 -1014
rect 138 -1028 146 -1027
rect 138 -1031 146 -1030
rect 172 -1083 180 -1082
rect 71 -1090 79 -1089
rect 172 -1086 180 -1085
rect 71 -1093 79 -1092
rect 71 -1115 79 -1114
rect 71 -1118 79 -1117
rect 172 -1119 180 -1118
rect 172 -1122 180 -1121
rect 71 -1140 79 -1139
rect 71 -1143 79 -1142
rect 172 -1144 180 -1143
rect 172 -1147 180 -1146
rect 172 -1169 180 -1168
rect 172 -1172 180 -1171
rect 59 -1185 67 -1184
rect 59 -1188 67 -1187
rect 172 -1194 180 -1193
rect 172 -1197 180 -1196
rect 59 -1210 67 -1209
rect 59 -1213 67 -1212
rect 172 -1219 180 -1218
rect 172 -1222 180 -1221
rect 59 -1235 67 -1234
rect 59 -1238 67 -1237
rect 303 -1441 311 -1440
rect 771 -1438 779 -1437
rect 532 -1441 540 -1440
rect -126 -1442 -118 -1441
rect -236 -1449 -228 -1448
rect -126 -1445 -118 -1444
rect 193 -1448 201 -1447
rect 303 -1444 311 -1443
rect 422 -1448 430 -1447
rect 532 -1444 540 -1443
rect 661 -1445 669 -1444
rect 771 -1441 779 -1440
rect -236 -1452 -228 -1451
rect 193 -1451 201 -1450
rect 422 -1451 430 -1450
rect 661 -1448 669 -1447
rect 193 -1473 201 -1472
rect -236 -1474 -228 -1473
rect -236 -1477 -228 -1476
rect -126 -1478 -118 -1477
rect 193 -1476 201 -1475
rect 661 -1470 669 -1469
rect 422 -1473 430 -1472
rect 303 -1477 311 -1476
rect -126 -1481 -118 -1480
rect 303 -1480 311 -1479
rect 422 -1476 430 -1475
rect 532 -1477 540 -1476
rect 661 -1473 669 -1472
rect 771 -1474 779 -1473
rect 532 -1480 540 -1479
rect 771 -1477 779 -1476
rect 193 -1498 201 -1497
rect -236 -1499 -228 -1498
rect -236 -1502 -228 -1501
rect -126 -1503 -118 -1502
rect 193 -1501 201 -1500
rect 661 -1495 669 -1494
rect 422 -1498 430 -1497
rect 303 -1502 311 -1501
rect -126 -1506 -118 -1505
rect 303 -1505 311 -1504
rect 422 -1501 430 -1500
rect 532 -1502 540 -1501
rect 661 -1498 669 -1497
rect 771 -1499 779 -1498
rect 532 -1505 540 -1504
rect 771 -1502 779 -1501
rect 303 -1527 311 -1526
rect 771 -1524 779 -1523
rect 532 -1527 540 -1526
rect -126 -1528 -118 -1527
rect -126 -1531 -118 -1530
rect 303 -1530 311 -1529
rect 532 -1530 540 -1529
rect 771 -1527 779 -1526
rect 303 -1552 311 -1551
rect 771 -1549 779 -1548
rect 532 -1552 540 -1551
rect -126 -1553 -118 -1552
rect -126 -1556 -118 -1555
rect 303 -1555 311 -1554
rect 532 -1555 540 -1554
rect 771 -1552 779 -1551
rect 303 -1577 311 -1576
rect 771 -1574 779 -1573
rect 532 -1577 540 -1576
rect -126 -1578 -118 -1577
rect -126 -1581 -118 -1580
rect 303 -1580 311 -1579
rect 532 -1580 540 -1579
rect 771 -1577 779 -1576
rect 337 -1632 345 -1631
rect 805 -1629 813 -1628
rect 566 -1632 574 -1631
rect -92 -1633 -84 -1632
rect -193 -1640 -185 -1639
rect -92 -1636 -84 -1635
rect 236 -1639 244 -1638
rect 337 -1635 345 -1634
rect 465 -1639 473 -1638
rect 566 -1635 574 -1634
rect 704 -1636 712 -1635
rect 805 -1632 813 -1631
rect -193 -1643 -185 -1642
rect 236 -1642 244 -1641
rect 465 -1642 473 -1641
rect 704 -1639 712 -1638
rect 236 -1664 244 -1663
rect -193 -1665 -185 -1664
rect -193 -1668 -185 -1667
rect -92 -1669 -84 -1668
rect 236 -1667 244 -1666
rect 704 -1661 712 -1660
rect 465 -1664 473 -1663
rect 337 -1668 345 -1667
rect -92 -1672 -84 -1671
rect 337 -1671 345 -1670
rect 465 -1667 473 -1666
rect 566 -1668 574 -1667
rect 704 -1664 712 -1663
rect 805 -1665 813 -1664
rect 566 -1671 574 -1670
rect 805 -1668 813 -1667
rect 236 -1689 244 -1688
rect -193 -1690 -185 -1689
rect -193 -1693 -185 -1692
rect -92 -1694 -84 -1693
rect 236 -1692 244 -1691
rect 704 -1686 712 -1685
rect 465 -1689 473 -1688
rect 337 -1693 345 -1692
rect -92 -1697 -84 -1696
rect 337 -1696 345 -1695
rect 465 -1692 473 -1691
rect 566 -1693 574 -1692
rect 704 -1689 712 -1688
rect 805 -1690 813 -1689
rect 566 -1696 574 -1695
rect 805 -1693 813 -1692
rect 337 -1718 345 -1717
rect 805 -1715 813 -1714
rect 566 -1718 574 -1717
rect -92 -1719 -84 -1718
rect -92 -1722 -84 -1721
rect 337 -1721 345 -1720
rect 566 -1721 574 -1720
rect 805 -1718 813 -1717
rect 224 -1734 232 -1733
rect 692 -1731 700 -1730
rect 453 -1734 461 -1733
rect -205 -1735 -197 -1734
rect -205 -1738 -197 -1737
rect 224 -1737 232 -1736
rect 453 -1737 461 -1736
rect 692 -1734 700 -1733
rect 337 -1743 345 -1742
rect 805 -1740 813 -1739
rect 566 -1743 574 -1742
rect -92 -1744 -84 -1743
rect -92 -1747 -84 -1746
rect 337 -1746 345 -1745
rect 566 -1746 574 -1745
rect 805 -1743 813 -1742
rect 224 -1759 232 -1758
rect 692 -1756 700 -1755
rect 453 -1759 461 -1758
rect -205 -1760 -197 -1759
rect -205 -1763 -197 -1762
rect 224 -1762 232 -1761
rect 453 -1762 461 -1761
rect 692 -1759 700 -1758
rect 337 -1768 345 -1767
rect 805 -1765 813 -1764
rect 566 -1768 574 -1767
rect -92 -1769 -84 -1768
rect -92 -1772 -84 -1771
rect 337 -1771 345 -1770
rect 566 -1771 574 -1770
rect 805 -1768 813 -1767
rect 224 -1784 232 -1783
rect 692 -1781 700 -1780
rect 453 -1784 461 -1783
rect -205 -1785 -197 -1784
rect -205 -1788 -197 -1787
rect 224 -1787 232 -1786
rect 453 -1787 461 -1786
rect 692 -1784 700 -1783
rect 553 -1909 561 -1908
rect 71 -1920 79 -1919
rect 443 -1916 451 -1915
rect 553 -1912 561 -1911
rect 746 -1917 754 -1916
rect 309 -1920 317 -1919
rect -39 -1927 -31 -1926
rect 71 -1923 79 -1922
rect 199 -1927 207 -1926
rect 309 -1923 317 -1922
rect 443 -1919 451 -1918
rect 636 -1924 644 -1923
rect 746 -1920 754 -1919
rect -39 -1930 -31 -1929
rect 199 -1930 207 -1929
rect 636 -1927 644 -1926
rect 443 -1941 451 -1940
rect -39 -1952 -31 -1951
rect -39 -1955 -31 -1954
rect 443 -1944 451 -1943
rect 553 -1945 561 -1944
rect 199 -1952 207 -1951
rect 71 -1956 79 -1955
rect 71 -1959 79 -1958
rect 199 -1955 207 -1954
rect 553 -1948 561 -1947
rect 636 -1949 644 -1948
rect 309 -1956 317 -1955
rect 636 -1952 644 -1951
rect 746 -1953 754 -1952
rect 309 -1959 317 -1958
rect 746 -1956 754 -1955
rect 443 -1966 451 -1965
rect -39 -1977 -31 -1976
rect -39 -1980 -31 -1979
rect 443 -1969 451 -1968
rect 553 -1970 561 -1969
rect 199 -1977 207 -1976
rect 71 -1981 79 -1980
rect 71 -1984 79 -1983
rect 199 -1980 207 -1979
rect 553 -1973 561 -1972
rect 636 -1974 644 -1973
rect 309 -1981 317 -1980
rect 636 -1977 644 -1976
rect 746 -1978 754 -1977
rect 309 -1984 317 -1983
rect 746 -1981 754 -1980
rect 553 -1995 561 -1994
rect 71 -2006 79 -2005
rect 553 -1998 561 -1997
rect 746 -2003 754 -2002
rect 309 -2006 317 -2005
rect 71 -2009 79 -2008
rect 309 -2009 317 -2008
rect 746 -2006 754 -2005
rect 553 -2020 561 -2019
rect 71 -2031 79 -2030
rect 553 -2023 561 -2022
rect 746 -2028 754 -2027
rect 309 -2031 317 -2030
rect 71 -2034 79 -2033
rect 309 -2034 317 -2033
rect 746 -2031 754 -2030
rect 553 -2045 561 -2044
rect 71 -2056 79 -2055
rect 553 -2048 561 -2047
rect 746 -2053 754 -2052
rect 309 -2056 317 -2055
rect 71 -2059 79 -2058
rect 309 -2059 317 -2058
rect 746 -2056 754 -2055
rect 105 -2111 113 -2110
rect 780 -2108 788 -2107
rect 343 -2111 351 -2110
rect 4 -2118 12 -2117
rect 105 -2114 113 -2113
rect 242 -2118 250 -2117
rect 343 -2114 351 -2113
rect 679 -2115 687 -2114
rect 780 -2111 788 -2110
rect 4 -2121 12 -2120
rect 242 -2121 250 -2120
rect 679 -2118 687 -2117
rect 4 -2143 12 -2142
rect 4 -2146 12 -2145
rect 679 -2140 687 -2139
rect 242 -2143 250 -2142
rect 105 -2147 113 -2146
rect 105 -2150 113 -2149
rect 242 -2146 250 -2145
rect 343 -2147 351 -2146
rect 679 -2143 687 -2142
rect 780 -2144 788 -2143
rect 343 -2150 351 -2149
rect 780 -2147 788 -2146
rect 4 -2168 12 -2167
rect 4 -2171 12 -2170
rect 679 -2165 687 -2164
rect 242 -2168 250 -2167
rect 105 -2172 113 -2171
rect 105 -2175 113 -2174
rect 242 -2171 250 -2170
rect 343 -2172 351 -2171
rect 679 -2168 687 -2167
rect 780 -2169 788 -2168
rect 343 -2175 351 -2174
rect 780 -2172 788 -2171
rect 105 -2197 113 -2196
rect 780 -2194 788 -2193
rect 343 -2197 351 -2196
rect 105 -2200 113 -2199
rect 343 -2200 351 -2199
rect 780 -2197 788 -2196
rect -8 -2213 0 -2212
rect 667 -2210 675 -2209
rect 230 -2213 238 -2212
rect -8 -2216 0 -2215
rect 230 -2216 238 -2215
rect 667 -2213 675 -2212
rect 105 -2222 113 -2221
rect 780 -2219 788 -2218
rect 343 -2222 351 -2221
rect 105 -2225 113 -2224
rect 343 -2225 351 -2224
rect 780 -2222 788 -2221
rect -8 -2238 0 -2237
rect 667 -2235 675 -2234
rect 230 -2238 238 -2237
rect -8 -2241 0 -2240
rect 230 -2241 238 -2240
rect 667 -2238 675 -2237
rect 105 -2247 113 -2246
rect 780 -2244 788 -2243
rect 343 -2247 351 -2246
rect 105 -2250 113 -2249
rect 343 -2250 351 -2249
rect 780 -2247 788 -2246
rect -8 -2263 0 -2262
rect 667 -2260 675 -2259
rect 230 -2263 238 -2262
rect -8 -2266 0 -2265
rect 230 -2266 238 -2265
rect 667 -2263 675 -2262
<< ndcontact >>
rect 20 -758 24 -754
rect 80 -758 84 -754
rect 140 -758 144 -754
rect 200 -758 204 -754
rect 260 -758 264 -754
rect 320 -758 324 -754
rect 380 -758 384 -754
rect 440 -758 444 -754
rect 500 -758 504 -754
rect 560 -758 564 -754
rect 620 -758 624 -754
rect 680 -758 684 -754
rect 740 -758 744 -754
rect 800 -758 804 -754
rect 860 -758 864 -754
rect 920 -758 924 -754
rect 20 -766 24 -762
rect 80 -766 84 -762
rect 140 -766 144 -762
rect 200 -766 204 -762
rect 260 -766 264 -762
rect 320 -766 324 -762
rect 380 -766 384 -762
rect 440 -766 444 -762
rect 500 -766 504 -762
rect 560 -766 564 -762
rect 620 -766 624 -762
rect 680 -766 684 -762
rect 740 -766 744 -762
rect 800 -766 804 -762
rect 860 -766 864 -762
rect 920 -766 924 -762
rect 20 -783 24 -779
rect 80 -783 84 -779
rect 140 -783 144 -779
rect 200 -783 204 -779
rect 260 -783 264 -779
rect 320 -783 324 -779
rect 380 -783 384 -779
rect 440 -783 444 -779
rect 500 -783 504 -779
rect 560 -783 564 -779
rect 620 -783 624 -779
rect 680 -783 684 -779
rect 740 -783 744 -779
rect 800 -783 804 -779
rect 860 -783 864 -779
rect 920 -783 924 -779
rect 20 -791 24 -787
rect 80 -791 84 -787
rect 140 -791 144 -787
rect 200 -791 204 -787
rect 260 -791 264 -787
rect 320 -791 324 -787
rect 380 -791 384 -787
rect 440 -791 444 -787
rect 500 -791 504 -787
rect 560 -791 564 -787
rect 620 -791 624 -787
rect 680 -791 684 -787
rect 740 -791 744 -787
rect 800 -791 804 -787
rect 860 -791 864 -787
rect 920 -791 924 -787
rect 20 -808 24 -804
rect 80 -808 84 -804
rect 140 -808 144 -804
rect 200 -808 204 -804
rect 260 -808 264 -804
rect 320 -808 324 -804
rect 380 -808 384 -804
rect 440 -808 444 -804
rect 500 -808 504 -804
rect 560 -808 564 -804
rect 620 -808 624 -804
rect 680 -808 684 -804
rect 740 -808 744 -804
rect 800 -808 804 -804
rect 860 -808 864 -804
rect 920 -808 924 -804
rect 20 -816 24 -812
rect 80 -816 84 -812
rect 140 -816 144 -812
rect 200 -816 204 -812
rect 260 -816 264 -812
rect 320 -816 324 -812
rect 380 -816 384 -812
rect 440 -816 444 -812
rect 500 -816 504 -812
rect 560 -816 564 -812
rect 620 -816 624 -812
rect 680 -816 684 -812
rect 740 -816 744 -812
rect 800 -816 804 -812
rect 860 -816 864 -812
rect 920 -816 924 -812
rect 416 -871 420 -867
rect 342 -878 346 -874
rect 416 -879 420 -875
rect 653 -875 657 -871
rect 836 -875 840 -871
rect 342 -886 346 -882
rect 579 -882 583 -878
rect 653 -883 657 -879
rect 762 -882 766 -878
rect 836 -883 840 -879
rect 71 -891 75 -887
rect 579 -890 583 -886
rect 762 -890 766 -886
rect -3 -898 1 -894
rect 71 -899 75 -895
rect -3 -906 1 -902
rect 342 -903 346 -899
rect 342 -911 346 -907
rect 452 -907 456 -903
rect 579 -907 583 -903
rect 762 -907 766 -903
rect 452 -915 456 -911
rect 579 -915 583 -911
rect 689 -911 693 -907
rect 689 -919 693 -915
rect 762 -915 766 -911
rect 872 -911 876 -907
rect 872 -919 876 -915
rect -3 -923 1 -919
rect -3 -931 1 -927
rect 107 -927 111 -923
rect 342 -928 346 -924
rect 107 -935 111 -931
rect 342 -936 346 -932
rect 416 -932 420 -928
rect 579 -932 583 -928
rect 762 -932 766 -928
rect 416 -940 420 -936
rect 579 -940 583 -936
rect 653 -936 657 -932
rect 653 -944 657 -940
rect 762 -940 766 -936
rect 836 -936 840 -932
rect 836 -944 840 -940
rect -3 -948 1 -944
rect -3 -956 1 -952
rect 71 -952 75 -948
rect 71 -960 75 -956
rect 416 -957 420 -953
rect 416 -965 420 -961
rect 653 -961 657 -957
rect 836 -961 840 -957
rect 653 -969 657 -965
rect 836 -969 840 -965
rect 71 -977 75 -973
rect 71 -985 75 -981
rect 452 -982 456 -978
rect 452 -990 456 -986
rect 689 -986 693 -982
rect 872 -986 876 -982
rect 689 -994 693 -990
rect 872 -994 876 -990
rect 107 -1002 111 -998
rect 107 -1010 111 -1006
rect 416 -1007 420 -1003
rect 416 -1015 420 -1011
rect 653 -1011 657 -1007
rect 836 -1011 840 -1007
rect 653 -1019 657 -1015
rect 836 -1019 840 -1015
rect 71 -1027 75 -1023
rect 71 -1035 75 -1031
rect 105 -1082 109 -1078
rect 40 -1089 44 -1085
rect 105 -1090 109 -1086
rect 40 -1097 44 -1093
rect 40 -1114 44 -1110
rect 40 -1122 44 -1118
rect 141 -1118 145 -1114
rect 141 -1126 145 -1122
rect 40 -1139 44 -1135
rect 40 -1147 44 -1143
rect 105 -1143 109 -1139
rect 105 -1151 109 -1147
rect 105 -1168 109 -1164
rect 105 -1176 109 -1172
rect 15 -1184 19 -1180
rect 15 -1192 19 -1188
rect 141 -1193 145 -1189
rect 141 -1201 145 -1197
rect 15 -1209 19 -1205
rect 15 -1217 19 -1213
rect 105 -1218 109 -1214
rect 105 -1226 109 -1222
rect 28 -1234 32 -1230
rect 28 -1242 32 -1238
rect -193 -1441 -189 -1437
rect 236 -1440 240 -1436
rect 465 -1440 469 -1436
rect 704 -1437 708 -1433
rect -267 -1448 -263 -1444
rect -193 -1449 -189 -1445
rect 162 -1447 166 -1443
rect 236 -1448 240 -1444
rect 391 -1447 395 -1443
rect 465 -1448 469 -1444
rect 630 -1444 634 -1440
rect 704 -1445 708 -1441
rect -267 -1456 -263 -1452
rect 162 -1455 166 -1451
rect 391 -1455 395 -1451
rect 630 -1452 634 -1448
rect -267 -1473 -263 -1469
rect 162 -1472 166 -1468
rect 391 -1472 395 -1468
rect -267 -1481 -263 -1477
rect -157 -1477 -153 -1473
rect 162 -1480 166 -1476
rect 272 -1476 276 -1472
rect 630 -1469 634 -1465
rect -157 -1485 -153 -1481
rect 272 -1484 276 -1480
rect 391 -1480 395 -1476
rect 501 -1476 505 -1472
rect 630 -1477 634 -1473
rect 740 -1473 744 -1469
rect 501 -1484 505 -1480
rect 740 -1481 744 -1477
rect -267 -1498 -263 -1494
rect 162 -1497 166 -1493
rect 391 -1497 395 -1493
rect -267 -1506 -263 -1502
rect -193 -1502 -189 -1498
rect 162 -1505 166 -1501
rect 236 -1501 240 -1497
rect 630 -1494 634 -1490
rect -193 -1510 -189 -1506
rect 236 -1509 240 -1505
rect 391 -1505 395 -1501
rect 465 -1501 469 -1497
rect 630 -1502 634 -1498
rect 704 -1498 708 -1494
rect 465 -1509 469 -1505
rect 704 -1506 708 -1502
rect -193 -1527 -189 -1523
rect 236 -1526 240 -1522
rect 465 -1526 469 -1522
rect 704 -1523 708 -1519
rect -193 -1535 -189 -1531
rect 236 -1534 240 -1530
rect 465 -1534 469 -1530
rect 704 -1531 708 -1527
rect -157 -1552 -153 -1548
rect 272 -1551 276 -1547
rect 501 -1551 505 -1547
rect 740 -1548 744 -1544
rect -157 -1560 -153 -1556
rect 272 -1559 276 -1555
rect 501 -1559 505 -1555
rect 740 -1556 744 -1552
rect -193 -1577 -189 -1573
rect 236 -1576 240 -1572
rect 465 -1576 469 -1572
rect 704 -1573 708 -1569
rect -193 -1585 -189 -1581
rect 236 -1584 240 -1580
rect 465 -1584 469 -1580
rect 704 -1581 708 -1577
rect -159 -1632 -155 -1628
rect 270 -1631 274 -1627
rect 499 -1631 503 -1627
rect 738 -1628 742 -1624
rect -224 -1639 -220 -1635
rect -159 -1640 -155 -1636
rect 205 -1638 209 -1634
rect 270 -1639 274 -1635
rect 434 -1638 438 -1634
rect 499 -1639 503 -1635
rect 673 -1635 677 -1631
rect 738 -1636 742 -1632
rect -224 -1647 -220 -1643
rect 205 -1646 209 -1642
rect 434 -1646 438 -1642
rect 673 -1643 677 -1639
rect -224 -1664 -220 -1660
rect 205 -1663 209 -1659
rect 434 -1663 438 -1659
rect -224 -1672 -220 -1668
rect -123 -1668 -119 -1664
rect 205 -1671 209 -1667
rect 306 -1667 310 -1663
rect 673 -1660 677 -1656
rect -123 -1676 -119 -1672
rect 306 -1675 310 -1671
rect 434 -1671 438 -1667
rect 535 -1667 539 -1663
rect 673 -1668 677 -1664
rect 774 -1664 778 -1660
rect 535 -1675 539 -1671
rect 774 -1672 778 -1668
rect -224 -1689 -220 -1685
rect 205 -1688 209 -1684
rect 434 -1688 438 -1684
rect -224 -1697 -220 -1693
rect -159 -1693 -155 -1689
rect 205 -1696 209 -1692
rect 270 -1692 274 -1688
rect 673 -1685 677 -1681
rect -159 -1701 -155 -1697
rect 270 -1700 274 -1696
rect 434 -1696 438 -1692
rect 499 -1692 503 -1688
rect 673 -1693 677 -1689
rect 738 -1689 742 -1685
rect 499 -1700 503 -1696
rect 738 -1697 742 -1693
rect -159 -1718 -155 -1714
rect 270 -1717 274 -1713
rect 499 -1717 503 -1713
rect 738 -1714 742 -1710
rect -159 -1726 -155 -1722
rect 270 -1725 274 -1721
rect 499 -1725 503 -1721
rect 738 -1722 742 -1718
rect -249 -1734 -245 -1730
rect 180 -1733 184 -1729
rect 409 -1733 413 -1729
rect 648 -1730 652 -1726
rect -249 -1742 -245 -1738
rect -123 -1743 -119 -1739
rect 180 -1741 184 -1737
rect 306 -1742 310 -1738
rect 409 -1741 413 -1737
rect 648 -1738 652 -1734
rect 535 -1742 539 -1738
rect 774 -1739 778 -1735
rect -123 -1751 -119 -1747
rect 306 -1750 310 -1746
rect 535 -1750 539 -1746
rect 774 -1747 778 -1743
rect -249 -1759 -245 -1755
rect 180 -1758 184 -1754
rect 409 -1758 413 -1754
rect 648 -1755 652 -1751
rect -249 -1767 -245 -1763
rect -159 -1768 -155 -1764
rect 180 -1766 184 -1762
rect 270 -1767 274 -1763
rect 409 -1766 413 -1762
rect 648 -1763 652 -1759
rect 499 -1767 503 -1763
rect 738 -1764 742 -1760
rect -159 -1776 -155 -1772
rect 270 -1775 274 -1771
rect 499 -1775 503 -1771
rect 738 -1772 742 -1768
rect -236 -1784 -232 -1780
rect 193 -1783 197 -1779
rect 422 -1783 426 -1779
rect 661 -1780 665 -1776
rect -236 -1792 -232 -1788
rect 193 -1791 197 -1787
rect 422 -1791 426 -1787
rect 661 -1788 665 -1784
rect 486 -1908 490 -1904
rect 412 -1915 416 -1911
rect 4 -1919 8 -1915
rect 242 -1919 246 -1915
rect 486 -1916 490 -1912
rect 679 -1916 683 -1912
rect -70 -1926 -66 -1922
rect 4 -1927 8 -1923
rect 168 -1926 172 -1922
rect 242 -1927 246 -1923
rect 412 -1923 416 -1919
rect 605 -1923 609 -1919
rect 679 -1924 683 -1920
rect -70 -1934 -66 -1930
rect 168 -1934 172 -1930
rect 605 -1931 609 -1927
rect 412 -1940 416 -1936
rect -70 -1951 -66 -1947
rect 168 -1951 172 -1947
rect -70 -1959 -66 -1955
rect 40 -1955 44 -1951
rect 412 -1948 416 -1944
rect 522 -1944 526 -1940
rect 40 -1963 44 -1959
rect 168 -1959 172 -1955
rect 278 -1955 282 -1951
rect 522 -1952 526 -1948
rect 605 -1948 609 -1944
rect 605 -1956 609 -1952
rect 715 -1952 719 -1948
rect 278 -1963 282 -1959
rect 715 -1960 719 -1956
rect 412 -1965 416 -1961
rect -70 -1976 -66 -1972
rect 168 -1976 172 -1972
rect -70 -1984 -66 -1980
rect 4 -1980 8 -1976
rect 412 -1973 416 -1969
rect 486 -1969 490 -1965
rect 4 -1988 8 -1984
rect 168 -1984 172 -1980
rect 242 -1980 246 -1976
rect 486 -1977 490 -1973
rect 605 -1973 609 -1969
rect 605 -1981 609 -1977
rect 679 -1977 683 -1973
rect 242 -1988 246 -1984
rect 679 -1985 683 -1981
rect 486 -1994 490 -1990
rect 4 -2005 8 -2001
rect 242 -2005 246 -2001
rect 486 -2002 490 -1998
rect 679 -2002 683 -1998
rect 4 -2013 8 -2009
rect 242 -2013 246 -2009
rect 679 -2010 683 -2006
rect 522 -2019 526 -2015
rect 40 -2030 44 -2026
rect 278 -2030 282 -2026
rect 522 -2027 526 -2023
rect 715 -2027 719 -2023
rect 40 -2038 44 -2034
rect 278 -2038 282 -2034
rect 715 -2035 719 -2031
rect 486 -2044 490 -2040
rect 4 -2055 8 -2051
rect 242 -2055 246 -2051
rect 486 -2052 490 -2048
rect 679 -2052 683 -2048
rect 4 -2063 8 -2059
rect 242 -2063 246 -2059
rect 679 -2060 683 -2056
rect 38 -2110 42 -2106
rect 276 -2110 280 -2106
rect 713 -2107 717 -2103
rect -27 -2117 -23 -2113
rect 38 -2118 42 -2114
rect 211 -2117 215 -2113
rect 276 -2118 280 -2114
rect 648 -2114 652 -2110
rect 713 -2115 717 -2111
rect -27 -2125 -23 -2121
rect 211 -2125 215 -2121
rect 648 -2122 652 -2118
rect -27 -2142 -23 -2138
rect 211 -2142 215 -2138
rect -27 -2150 -23 -2146
rect 74 -2146 78 -2142
rect 648 -2139 652 -2135
rect 74 -2154 78 -2150
rect 211 -2150 215 -2146
rect 312 -2146 316 -2142
rect 648 -2147 652 -2143
rect 749 -2143 753 -2139
rect 312 -2154 316 -2150
rect 749 -2151 753 -2147
rect -27 -2167 -23 -2163
rect 211 -2167 215 -2163
rect -27 -2175 -23 -2171
rect 38 -2171 42 -2167
rect 648 -2164 652 -2160
rect 38 -2179 42 -2175
rect 211 -2175 215 -2171
rect 276 -2171 280 -2167
rect 648 -2172 652 -2168
rect 713 -2168 717 -2164
rect 276 -2179 280 -2175
rect 713 -2176 717 -2172
rect 38 -2196 42 -2192
rect 276 -2196 280 -2192
rect 713 -2193 717 -2189
rect 38 -2204 42 -2200
rect 276 -2204 280 -2200
rect 713 -2201 717 -2197
rect -52 -2212 -48 -2208
rect 186 -2212 190 -2208
rect 623 -2209 627 -2205
rect -52 -2220 -48 -2216
rect 74 -2221 78 -2217
rect 186 -2220 190 -2216
rect 623 -2217 627 -2213
rect 312 -2221 316 -2217
rect 749 -2218 753 -2214
rect 74 -2229 78 -2225
rect 312 -2229 316 -2225
rect 749 -2226 753 -2222
rect -52 -2237 -48 -2233
rect 186 -2237 190 -2233
rect 623 -2234 627 -2230
rect -52 -2245 -48 -2241
rect 38 -2246 42 -2242
rect 186 -2245 190 -2241
rect 623 -2242 627 -2238
rect 276 -2246 280 -2242
rect 713 -2243 717 -2239
rect 38 -2254 42 -2250
rect 276 -2254 280 -2250
rect 713 -2251 717 -2247
rect -39 -2262 -35 -2258
rect 199 -2262 203 -2258
rect 636 -2259 640 -2255
rect -39 -2270 -35 -2266
rect 199 -2270 203 -2266
rect 636 -2267 640 -2263
<< pdcontact >>
rect 51 -758 59 -754
rect 111 -758 119 -754
rect 171 -758 179 -754
rect 231 -758 239 -754
rect 291 -758 299 -754
rect 351 -758 359 -754
rect 411 -758 419 -754
rect 471 -758 479 -754
rect 531 -758 539 -754
rect 591 -758 599 -754
rect 651 -758 659 -754
rect 711 -758 719 -754
rect 771 -758 779 -754
rect 831 -758 839 -754
rect 891 -758 899 -754
rect 951 -758 959 -754
rect 51 -766 59 -762
rect 111 -766 119 -762
rect 171 -766 179 -762
rect 231 -766 239 -762
rect 291 -766 299 -762
rect 351 -766 359 -762
rect 411 -766 419 -762
rect 471 -766 479 -762
rect 531 -766 539 -762
rect 591 -766 599 -762
rect 651 -766 659 -762
rect 711 -766 719 -762
rect 771 -766 779 -762
rect 831 -766 839 -762
rect 891 -766 899 -762
rect 951 -766 959 -762
rect 51 -783 59 -779
rect 111 -783 119 -779
rect 171 -783 179 -779
rect 231 -783 239 -779
rect 291 -783 299 -779
rect 351 -783 359 -779
rect 411 -783 419 -779
rect 471 -783 479 -779
rect 531 -783 539 -779
rect 591 -783 599 -779
rect 651 -783 659 -779
rect 711 -783 719 -779
rect 771 -783 779 -779
rect 831 -783 839 -779
rect 891 -783 899 -779
rect 951 -783 959 -779
rect 51 -791 59 -787
rect 111 -791 119 -787
rect 171 -791 179 -787
rect 231 -791 239 -787
rect 291 -791 299 -787
rect 351 -791 359 -787
rect 411 -791 419 -787
rect 471 -791 479 -787
rect 531 -791 539 -787
rect 591 -791 599 -787
rect 651 -791 659 -787
rect 711 -791 719 -787
rect 771 -791 779 -787
rect 831 -791 839 -787
rect 891 -791 899 -787
rect 951 -791 959 -787
rect 51 -808 59 -804
rect 111 -808 119 -804
rect 171 -808 179 -804
rect 231 -808 239 -804
rect 291 -808 299 -804
rect 351 -808 359 -804
rect 411 -808 419 -804
rect 471 -808 479 -804
rect 531 -808 539 -804
rect 591 -808 599 -804
rect 651 -808 659 -804
rect 711 -808 719 -804
rect 771 -808 779 -804
rect 831 -808 839 -804
rect 891 -808 899 -804
rect 951 -808 959 -804
rect 51 -816 59 -812
rect 111 -816 119 -812
rect 171 -816 179 -812
rect 231 -816 239 -812
rect 291 -816 299 -812
rect 351 -816 359 -812
rect 411 -816 419 -812
rect 471 -816 479 -812
rect 531 -816 539 -812
rect 591 -816 599 -812
rect 651 -816 659 -812
rect 711 -816 719 -812
rect 771 -816 779 -812
rect 831 -816 839 -812
rect 891 -816 899 -812
rect 951 -816 959 -812
rect 483 -871 491 -867
rect 373 -878 381 -874
rect 483 -879 491 -875
rect 720 -875 728 -871
rect 903 -875 911 -871
rect 373 -886 381 -882
rect 610 -882 618 -878
rect 720 -883 728 -879
rect 793 -882 801 -878
rect 903 -883 911 -879
rect 138 -891 146 -887
rect 610 -890 618 -886
rect 793 -890 801 -886
rect 28 -898 36 -894
rect 138 -899 146 -895
rect 28 -906 36 -902
rect 373 -903 381 -899
rect 373 -911 381 -907
rect 483 -907 491 -903
rect 610 -907 618 -903
rect 483 -915 491 -911
rect 610 -915 618 -911
rect 720 -911 728 -907
rect 793 -907 801 -903
rect 793 -915 801 -911
rect 903 -911 911 -907
rect 720 -919 728 -915
rect 903 -919 911 -915
rect 28 -923 36 -919
rect 28 -931 36 -927
rect 138 -927 146 -923
rect 373 -928 381 -924
rect 138 -935 146 -931
rect 373 -936 381 -932
rect 483 -932 491 -928
rect 610 -932 618 -928
rect 483 -940 491 -936
rect 610 -940 618 -936
rect 720 -936 728 -932
rect 793 -932 801 -928
rect 793 -940 801 -936
rect 903 -936 911 -932
rect 720 -944 728 -940
rect 903 -944 911 -940
rect 28 -948 36 -944
rect 28 -956 36 -952
rect 138 -952 146 -948
rect 138 -960 146 -956
rect 483 -957 491 -953
rect 483 -965 491 -961
rect 720 -961 728 -957
rect 903 -961 911 -957
rect 720 -969 728 -965
rect 903 -969 911 -965
rect 138 -977 146 -973
rect 138 -985 146 -981
rect 483 -982 491 -978
rect 483 -990 491 -986
rect 720 -986 728 -982
rect 903 -986 911 -982
rect 720 -994 728 -990
rect 903 -994 911 -990
rect 138 -1002 146 -998
rect 138 -1010 146 -1006
rect 483 -1007 491 -1003
rect 483 -1015 491 -1011
rect 720 -1011 728 -1007
rect 903 -1011 911 -1007
rect 720 -1019 728 -1015
rect 903 -1019 911 -1015
rect 138 -1027 146 -1023
rect 138 -1035 146 -1031
rect 172 -1082 180 -1078
rect 71 -1089 79 -1085
rect 172 -1090 180 -1086
rect 71 -1097 79 -1093
rect 71 -1114 79 -1110
rect 71 -1122 79 -1118
rect 172 -1118 180 -1114
rect 172 -1126 180 -1122
rect 71 -1139 79 -1135
rect 71 -1147 79 -1143
rect 172 -1143 180 -1139
rect 172 -1151 180 -1147
rect 172 -1168 180 -1164
rect 172 -1176 180 -1172
rect 59 -1184 67 -1180
rect 59 -1192 67 -1188
rect 172 -1193 180 -1189
rect 172 -1201 180 -1197
rect 59 -1209 67 -1205
rect 59 -1217 67 -1213
rect 172 -1218 180 -1214
rect 172 -1226 180 -1222
rect 59 -1234 67 -1230
rect 59 -1242 67 -1238
rect -126 -1441 -118 -1437
rect 303 -1440 311 -1436
rect 532 -1440 540 -1436
rect 771 -1437 779 -1433
rect -236 -1448 -228 -1444
rect -126 -1449 -118 -1445
rect 193 -1447 201 -1443
rect 303 -1448 311 -1444
rect 422 -1447 430 -1443
rect 532 -1448 540 -1444
rect 661 -1444 669 -1440
rect 771 -1445 779 -1441
rect -236 -1456 -228 -1452
rect 193 -1455 201 -1451
rect 422 -1455 430 -1451
rect 661 -1452 669 -1448
rect -236 -1473 -228 -1469
rect 193 -1472 201 -1468
rect -236 -1481 -228 -1477
rect -126 -1477 -118 -1473
rect 193 -1480 201 -1476
rect 303 -1476 311 -1472
rect 422 -1472 430 -1468
rect 661 -1469 669 -1465
rect -126 -1485 -118 -1481
rect 422 -1480 430 -1476
rect 532 -1476 540 -1472
rect 661 -1477 669 -1473
rect 771 -1473 779 -1469
rect 303 -1484 311 -1480
rect 532 -1484 540 -1480
rect 771 -1481 779 -1477
rect -236 -1498 -228 -1494
rect 193 -1497 201 -1493
rect -236 -1506 -228 -1502
rect -126 -1502 -118 -1498
rect 193 -1505 201 -1501
rect 303 -1501 311 -1497
rect 422 -1497 430 -1493
rect 661 -1494 669 -1490
rect -126 -1510 -118 -1506
rect 422 -1505 430 -1501
rect 532 -1501 540 -1497
rect 661 -1502 669 -1498
rect 771 -1498 779 -1494
rect 303 -1509 311 -1505
rect 532 -1509 540 -1505
rect 771 -1506 779 -1502
rect -126 -1527 -118 -1523
rect 303 -1526 311 -1522
rect 532 -1526 540 -1522
rect 771 -1523 779 -1519
rect -126 -1535 -118 -1531
rect 303 -1534 311 -1530
rect 532 -1534 540 -1530
rect 771 -1531 779 -1527
rect -126 -1552 -118 -1548
rect 303 -1551 311 -1547
rect 532 -1551 540 -1547
rect 771 -1548 779 -1544
rect -126 -1560 -118 -1556
rect 303 -1559 311 -1555
rect 532 -1559 540 -1555
rect 771 -1556 779 -1552
rect -126 -1577 -118 -1573
rect 303 -1576 311 -1572
rect 532 -1576 540 -1572
rect 771 -1573 779 -1569
rect -126 -1585 -118 -1581
rect 303 -1584 311 -1580
rect 532 -1584 540 -1580
rect 771 -1581 779 -1577
rect -92 -1632 -84 -1628
rect 337 -1631 345 -1627
rect 566 -1631 574 -1627
rect 805 -1628 813 -1624
rect -193 -1639 -185 -1635
rect -92 -1640 -84 -1636
rect 236 -1638 244 -1634
rect 337 -1639 345 -1635
rect 465 -1638 473 -1634
rect 566 -1639 574 -1635
rect 704 -1635 712 -1631
rect 805 -1636 813 -1632
rect -193 -1647 -185 -1643
rect 236 -1646 244 -1642
rect 465 -1646 473 -1642
rect 704 -1643 712 -1639
rect -193 -1664 -185 -1660
rect 236 -1663 244 -1659
rect -193 -1672 -185 -1668
rect -92 -1668 -84 -1664
rect 236 -1671 244 -1667
rect 337 -1667 345 -1663
rect 465 -1663 473 -1659
rect 704 -1660 712 -1656
rect -92 -1676 -84 -1672
rect 465 -1671 473 -1667
rect 566 -1667 574 -1663
rect 704 -1668 712 -1664
rect 805 -1664 813 -1660
rect 337 -1675 345 -1671
rect 566 -1675 574 -1671
rect 805 -1672 813 -1668
rect -193 -1689 -185 -1685
rect 236 -1688 244 -1684
rect -193 -1697 -185 -1693
rect -92 -1693 -84 -1689
rect 236 -1696 244 -1692
rect 337 -1692 345 -1688
rect 465 -1688 473 -1684
rect 704 -1685 712 -1681
rect -92 -1701 -84 -1697
rect 465 -1696 473 -1692
rect 566 -1692 574 -1688
rect 704 -1693 712 -1689
rect 805 -1689 813 -1685
rect 337 -1700 345 -1696
rect 566 -1700 574 -1696
rect 805 -1697 813 -1693
rect -92 -1718 -84 -1714
rect 337 -1717 345 -1713
rect 566 -1717 574 -1713
rect 805 -1714 813 -1710
rect -92 -1726 -84 -1722
rect 337 -1725 345 -1721
rect 566 -1725 574 -1721
rect 805 -1722 813 -1718
rect -205 -1734 -197 -1730
rect 224 -1733 232 -1729
rect 453 -1733 461 -1729
rect 692 -1730 700 -1726
rect -205 -1742 -197 -1738
rect -92 -1743 -84 -1739
rect 224 -1741 232 -1737
rect 337 -1742 345 -1738
rect 453 -1741 461 -1737
rect 692 -1738 700 -1734
rect 566 -1742 574 -1738
rect 805 -1739 813 -1735
rect -92 -1751 -84 -1747
rect 337 -1750 345 -1746
rect 566 -1750 574 -1746
rect 805 -1747 813 -1743
rect -205 -1759 -197 -1755
rect 224 -1758 232 -1754
rect 453 -1758 461 -1754
rect 692 -1755 700 -1751
rect -205 -1767 -197 -1763
rect -92 -1768 -84 -1764
rect 224 -1766 232 -1762
rect 337 -1767 345 -1763
rect 453 -1766 461 -1762
rect 692 -1763 700 -1759
rect 566 -1767 574 -1763
rect 805 -1764 813 -1760
rect -92 -1776 -84 -1772
rect 337 -1775 345 -1771
rect 566 -1775 574 -1771
rect 805 -1772 813 -1768
rect -205 -1784 -197 -1780
rect 224 -1783 232 -1779
rect 453 -1783 461 -1779
rect 692 -1780 700 -1776
rect -205 -1792 -197 -1788
rect 224 -1791 232 -1787
rect 453 -1791 461 -1787
rect 692 -1788 700 -1784
rect 553 -1908 561 -1904
rect 71 -1919 79 -1915
rect 309 -1919 317 -1915
rect 443 -1915 451 -1911
rect 553 -1916 561 -1912
rect 746 -1916 754 -1912
rect -39 -1926 -31 -1922
rect 71 -1927 79 -1923
rect 199 -1926 207 -1922
rect 443 -1923 451 -1919
rect 309 -1927 317 -1923
rect 636 -1923 644 -1919
rect 746 -1924 754 -1920
rect -39 -1934 -31 -1930
rect 199 -1934 207 -1930
rect 636 -1931 644 -1927
rect 443 -1940 451 -1936
rect -39 -1951 -31 -1947
rect -39 -1959 -31 -1955
rect 71 -1955 79 -1951
rect 199 -1951 207 -1947
rect 443 -1948 451 -1944
rect 553 -1944 561 -1940
rect 199 -1959 207 -1955
rect 309 -1955 317 -1951
rect 553 -1952 561 -1948
rect 636 -1948 644 -1944
rect 636 -1956 644 -1952
rect 746 -1952 754 -1948
rect 71 -1963 79 -1959
rect 309 -1963 317 -1959
rect 746 -1960 754 -1956
rect 443 -1965 451 -1961
rect -39 -1976 -31 -1972
rect -39 -1984 -31 -1980
rect 71 -1980 79 -1976
rect 199 -1976 207 -1972
rect 443 -1973 451 -1969
rect 553 -1969 561 -1965
rect 199 -1984 207 -1980
rect 309 -1980 317 -1976
rect 553 -1977 561 -1973
rect 636 -1973 644 -1969
rect 636 -1981 644 -1977
rect 746 -1977 754 -1973
rect 71 -1988 79 -1984
rect 309 -1988 317 -1984
rect 746 -1985 754 -1981
rect 553 -1994 561 -1990
rect 71 -2005 79 -2001
rect 309 -2005 317 -2001
rect 553 -2002 561 -1998
rect 746 -2002 754 -1998
rect 71 -2013 79 -2009
rect 309 -2013 317 -2009
rect 746 -2010 754 -2006
rect 553 -2019 561 -2015
rect 71 -2030 79 -2026
rect 309 -2030 317 -2026
rect 553 -2027 561 -2023
rect 746 -2027 754 -2023
rect 71 -2038 79 -2034
rect 309 -2038 317 -2034
rect 746 -2035 754 -2031
rect 553 -2044 561 -2040
rect 71 -2055 79 -2051
rect 309 -2055 317 -2051
rect 553 -2052 561 -2048
rect 746 -2052 754 -2048
rect 71 -2063 79 -2059
rect 309 -2063 317 -2059
rect 746 -2060 754 -2056
rect 105 -2110 113 -2106
rect 343 -2110 351 -2106
rect 780 -2107 788 -2103
rect 4 -2117 12 -2113
rect 105 -2118 113 -2114
rect 242 -2117 250 -2113
rect 343 -2118 351 -2114
rect 679 -2114 687 -2110
rect 780 -2115 788 -2111
rect 4 -2125 12 -2121
rect 242 -2125 250 -2121
rect 679 -2122 687 -2118
rect 4 -2142 12 -2138
rect 4 -2150 12 -2146
rect 105 -2146 113 -2142
rect 242 -2142 250 -2138
rect 679 -2139 687 -2135
rect 242 -2150 250 -2146
rect 343 -2146 351 -2142
rect 679 -2147 687 -2143
rect 780 -2143 788 -2139
rect 105 -2154 113 -2150
rect 343 -2154 351 -2150
rect 780 -2151 788 -2147
rect 4 -2167 12 -2163
rect 4 -2175 12 -2171
rect 105 -2171 113 -2167
rect 242 -2167 250 -2163
rect 679 -2164 687 -2160
rect 242 -2175 250 -2171
rect 343 -2171 351 -2167
rect 679 -2172 687 -2168
rect 780 -2168 788 -2164
rect 105 -2179 113 -2175
rect 343 -2179 351 -2175
rect 780 -2176 788 -2172
rect 105 -2196 113 -2192
rect 343 -2196 351 -2192
rect 780 -2193 788 -2189
rect 105 -2204 113 -2200
rect 343 -2204 351 -2200
rect 780 -2201 788 -2197
rect -8 -2212 0 -2208
rect 230 -2212 238 -2208
rect 667 -2209 675 -2205
rect -8 -2220 0 -2216
rect 105 -2221 113 -2217
rect 230 -2220 238 -2216
rect 667 -2217 675 -2213
rect 343 -2221 351 -2217
rect 780 -2218 788 -2214
rect 105 -2229 113 -2225
rect 343 -2229 351 -2225
rect 780 -2226 788 -2222
rect -8 -2237 0 -2233
rect 230 -2237 238 -2233
rect 667 -2234 675 -2230
rect -8 -2245 0 -2241
rect 105 -2246 113 -2242
rect 230 -2245 238 -2241
rect 667 -2242 675 -2238
rect 343 -2246 351 -2242
rect 780 -2243 788 -2239
rect 105 -2254 113 -2250
rect 343 -2254 351 -2250
rect 780 -2251 788 -2247
rect -8 -2262 0 -2258
rect 230 -2262 238 -2258
rect 667 -2259 675 -2255
rect -8 -2270 0 -2266
rect 230 -2270 238 -2266
rect 667 -2267 675 -2263
<< polysilicon >>
rect 17 -761 20 -759
rect 24 -761 51 -759
rect 59 -761 62 -759
rect 77 -761 80 -759
rect 84 -761 111 -759
rect 119 -761 122 -759
rect 137 -761 140 -759
rect 144 -761 171 -759
rect 179 -761 182 -759
rect 197 -761 200 -759
rect 204 -761 231 -759
rect 239 -761 242 -759
rect 257 -761 260 -759
rect 264 -761 291 -759
rect 299 -761 302 -759
rect 317 -761 320 -759
rect 324 -761 351 -759
rect 359 -761 362 -759
rect 377 -761 380 -759
rect 384 -761 411 -759
rect 419 -761 422 -759
rect 437 -761 440 -759
rect 444 -761 471 -759
rect 479 -761 482 -759
rect 497 -761 500 -759
rect 504 -761 531 -759
rect 539 -761 542 -759
rect 557 -761 560 -759
rect 564 -761 591 -759
rect 599 -761 602 -759
rect 617 -761 620 -759
rect 624 -761 651 -759
rect 659 -761 662 -759
rect 677 -761 680 -759
rect 684 -761 711 -759
rect 719 -761 722 -759
rect 737 -761 740 -759
rect 744 -761 771 -759
rect 779 -761 782 -759
rect 797 -761 800 -759
rect 804 -761 831 -759
rect 839 -761 842 -759
rect 857 -761 860 -759
rect 864 -761 891 -759
rect 899 -761 902 -759
rect 917 -761 920 -759
rect 924 -761 951 -759
rect 959 -761 962 -759
rect 17 -786 20 -784
rect 24 -786 51 -784
rect 59 -786 62 -784
rect 77 -786 80 -784
rect 84 -786 111 -784
rect 119 -786 122 -784
rect 137 -786 140 -784
rect 144 -786 171 -784
rect 179 -786 182 -784
rect 197 -786 200 -784
rect 204 -786 231 -784
rect 239 -786 242 -784
rect 257 -786 260 -784
rect 264 -786 291 -784
rect 299 -786 302 -784
rect 317 -786 320 -784
rect 324 -786 351 -784
rect 359 -786 362 -784
rect 377 -786 380 -784
rect 384 -786 411 -784
rect 419 -786 422 -784
rect 437 -786 440 -784
rect 444 -786 471 -784
rect 479 -786 482 -784
rect 497 -786 500 -784
rect 504 -786 531 -784
rect 539 -786 542 -784
rect 557 -786 560 -784
rect 564 -786 591 -784
rect 599 -786 602 -784
rect 617 -786 620 -784
rect 624 -786 651 -784
rect 659 -786 662 -784
rect 677 -786 680 -784
rect 684 -786 711 -784
rect 719 -786 722 -784
rect 737 -786 740 -784
rect 744 -786 771 -784
rect 779 -786 782 -784
rect 797 -786 800 -784
rect 804 -786 831 -784
rect 839 -786 842 -784
rect 857 -786 860 -784
rect 864 -786 891 -784
rect 899 -786 902 -784
rect 917 -786 920 -784
rect 924 -786 951 -784
rect 959 -786 962 -784
rect 17 -811 20 -809
rect 24 -811 51 -809
rect 59 -811 62 -809
rect 77 -811 80 -809
rect 84 -811 111 -809
rect 119 -811 122 -809
rect 137 -811 140 -809
rect 144 -811 171 -809
rect 179 -811 182 -809
rect 197 -811 200 -809
rect 204 -811 231 -809
rect 239 -811 242 -809
rect 257 -811 260 -809
rect 264 -811 291 -809
rect 299 -811 302 -809
rect 317 -811 320 -809
rect 324 -811 351 -809
rect 359 -811 362 -809
rect 377 -811 380 -809
rect 384 -811 411 -809
rect 419 -811 422 -809
rect 437 -811 440 -809
rect 444 -811 471 -809
rect 479 -811 482 -809
rect 497 -811 500 -809
rect 504 -811 531 -809
rect 539 -811 542 -809
rect 557 -811 560 -809
rect 564 -811 591 -809
rect 599 -811 602 -809
rect 617 -811 620 -809
rect 624 -811 651 -809
rect 659 -811 662 -809
rect 677 -811 680 -809
rect 684 -811 711 -809
rect 719 -811 722 -809
rect 737 -811 740 -809
rect 744 -811 771 -809
rect 779 -811 782 -809
rect 797 -811 800 -809
rect 804 -811 831 -809
rect 839 -811 842 -809
rect 857 -811 860 -809
rect 864 -811 891 -809
rect 899 -811 902 -809
rect 917 -811 920 -809
rect 924 -811 951 -809
rect 959 -811 962 -809
rect 413 -874 416 -872
rect 420 -874 483 -872
rect 491 -874 494 -872
rect 650 -878 653 -876
rect 657 -878 720 -876
rect 728 -878 731 -876
rect 833 -878 836 -876
rect 840 -878 903 -876
rect 911 -878 914 -876
rect 339 -881 342 -879
rect 346 -881 373 -879
rect 381 -881 384 -879
rect 576 -885 579 -883
rect 583 -885 610 -883
rect 618 -885 621 -883
rect 759 -885 762 -883
rect 766 -885 793 -883
rect 801 -885 804 -883
rect 68 -894 71 -892
rect 75 -894 138 -892
rect 146 -894 149 -892
rect -6 -901 -3 -899
rect 1 -901 28 -899
rect 36 -901 39 -899
rect 339 -906 342 -904
rect 346 -906 373 -904
rect 381 -906 384 -904
rect 449 -910 452 -908
rect 456 -910 483 -908
rect 491 -910 494 -908
rect 576 -910 579 -908
rect 583 -910 610 -908
rect 618 -910 621 -908
rect 759 -910 762 -908
rect 766 -910 793 -908
rect 801 -910 804 -908
rect 686 -914 689 -912
rect 693 -914 720 -912
rect 728 -914 731 -912
rect 869 -914 872 -912
rect 876 -914 903 -912
rect 911 -914 914 -912
rect -6 -926 -3 -924
rect 1 -926 28 -924
rect 36 -926 39 -924
rect 104 -930 107 -928
rect 111 -930 138 -928
rect 146 -930 149 -928
rect 339 -931 342 -929
rect 346 -931 373 -929
rect 381 -931 384 -929
rect 413 -935 416 -933
rect 420 -935 483 -933
rect 491 -935 494 -933
rect 576 -935 579 -933
rect 583 -935 610 -933
rect 618 -935 621 -933
rect 759 -935 762 -933
rect 766 -935 793 -933
rect 801 -935 804 -933
rect 650 -939 653 -937
rect 657 -939 720 -937
rect 728 -939 731 -937
rect 833 -939 836 -937
rect 840 -939 903 -937
rect 911 -939 914 -937
rect -6 -951 -3 -949
rect 1 -951 28 -949
rect 36 -951 39 -949
rect 68 -955 71 -953
rect 75 -955 138 -953
rect 146 -955 149 -953
rect 413 -960 416 -958
rect 420 -960 483 -958
rect 491 -960 494 -958
rect 650 -964 653 -962
rect 657 -964 720 -962
rect 728 -964 731 -962
rect 833 -964 836 -962
rect 840 -964 903 -962
rect 911 -964 914 -962
rect 68 -980 71 -978
rect 75 -980 138 -978
rect 146 -980 149 -978
rect 449 -985 452 -983
rect 456 -985 483 -983
rect 491 -985 494 -983
rect 686 -989 689 -987
rect 693 -989 720 -987
rect 728 -989 731 -987
rect 869 -989 872 -987
rect 876 -989 903 -987
rect 911 -989 914 -987
rect 104 -1005 107 -1003
rect 111 -1005 138 -1003
rect 146 -1005 149 -1003
rect 413 -1010 416 -1008
rect 420 -1010 483 -1008
rect 491 -1010 494 -1008
rect 650 -1014 653 -1012
rect 657 -1014 720 -1012
rect 728 -1014 731 -1012
rect 833 -1014 836 -1012
rect 840 -1014 903 -1012
rect 911 -1014 914 -1012
rect 68 -1030 71 -1028
rect 75 -1030 138 -1028
rect 146 -1030 149 -1028
rect 102 -1085 105 -1083
rect 109 -1085 172 -1083
rect 180 -1085 183 -1083
rect 37 -1092 40 -1090
rect 44 -1092 71 -1090
rect 79 -1092 82 -1090
rect 37 -1117 40 -1115
rect 44 -1117 71 -1115
rect 79 -1117 82 -1115
rect 138 -1121 141 -1119
rect 145 -1121 172 -1119
rect 180 -1121 183 -1119
rect 37 -1142 40 -1140
rect 44 -1142 71 -1140
rect 79 -1142 82 -1140
rect 102 -1146 105 -1144
rect 109 -1146 172 -1144
rect 180 -1146 183 -1144
rect 102 -1171 105 -1169
rect 109 -1171 172 -1169
rect 180 -1171 183 -1169
rect 12 -1187 15 -1185
rect 19 -1187 59 -1185
rect 67 -1187 70 -1185
rect 138 -1196 141 -1194
rect 145 -1196 172 -1194
rect 180 -1196 183 -1194
rect 12 -1212 15 -1210
rect 19 -1212 59 -1210
rect 67 -1212 70 -1210
rect 102 -1221 105 -1219
rect 109 -1221 172 -1219
rect 180 -1221 183 -1219
rect 25 -1237 28 -1235
rect 32 -1237 59 -1235
rect 67 -1237 70 -1235
rect 701 -1440 704 -1438
rect 708 -1440 771 -1438
rect 779 -1440 782 -1438
rect -196 -1444 -193 -1442
rect -189 -1444 -126 -1442
rect -118 -1444 -115 -1442
rect 233 -1443 236 -1441
rect 240 -1443 303 -1441
rect 311 -1443 314 -1441
rect 462 -1443 465 -1441
rect 469 -1443 532 -1441
rect 540 -1443 543 -1441
rect 627 -1447 630 -1445
rect 634 -1447 661 -1445
rect 669 -1447 672 -1445
rect -270 -1451 -267 -1449
rect -263 -1451 -236 -1449
rect -228 -1451 -225 -1449
rect 159 -1450 162 -1448
rect 166 -1450 193 -1448
rect 201 -1450 204 -1448
rect 388 -1450 391 -1448
rect 395 -1450 422 -1448
rect 430 -1450 433 -1448
rect -270 -1476 -267 -1474
rect -263 -1476 -236 -1474
rect -228 -1476 -225 -1474
rect 159 -1475 162 -1473
rect 166 -1475 193 -1473
rect 201 -1475 204 -1473
rect -160 -1480 -157 -1478
rect -153 -1480 -126 -1478
rect -118 -1480 -115 -1478
rect 627 -1472 630 -1470
rect 634 -1472 661 -1470
rect 669 -1472 672 -1470
rect 388 -1475 391 -1473
rect 395 -1475 422 -1473
rect 430 -1475 433 -1473
rect 269 -1479 272 -1477
rect 276 -1479 303 -1477
rect 311 -1479 314 -1477
rect 737 -1476 740 -1474
rect 744 -1476 771 -1474
rect 779 -1476 782 -1474
rect 498 -1479 501 -1477
rect 505 -1479 532 -1477
rect 540 -1479 543 -1477
rect -270 -1501 -267 -1499
rect -263 -1501 -236 -1499
rect -228 -1501 -225 -1499
rect 159 -1500 162 -1498
rect 166 -1500 193 -1498
rect 201 -1500 204 -1498
rect -196 -1505 -193 -1503
rect -189 -1505 -126 -1503
rect -118 -1505 -115 -1503
rect 627 -1497 630 -1495
rect 634 -1497 661 -1495
rect 669 -1497 672 -1495
rect 388 -1500 391 -1498
rect 395 -1500 422 -1498
rect 430 -1500 433 -1498
rect 233 -1504 236 -1502
rect 240 -1504 303 -1502
rect 311 -1504 314 -1502
rect 701 -1501 704 -1499
rect 708 -1501 771 -1499
rect 779 -1501 782 -1499
rect 462 -1504 465 -1502
rect 469 -1504 532 -1502
rect 540 -1504 543 -1502
rect 701 -1526 704 -1524
rect 708 -1526 771 -1524
rect 779 -1526 782 -1524
rect -196 -1530 -193 -1528
rect -189 -1530 -126 -1528
rect -118 -1530 -115 -1528
rect 233 -1529 236 -1527
rect 240 -1529 303 -1527
rect 311 -1529 314 -1527
rect 462 -1529 465 -1527
rect 469 -1529 532 -1527
rect 540 -1529 543 -1527
rect 737 -1551 740 -1549
rect 744 -1551 771 -1549
rect 779 -1551 782 -1549
rect -160 -1555 -157 -1553
rect -153 -1555 -126 -1553
rect -118 -1555 -115 -1553
rect 269 -1554 272 -1552
rect 276 -1554 303 -1552
rect 311 -1554 314 -1552
rect 498 -1554 501 -1552
rect 505 -1554 532 -1552
rect 540 -1554 543 -1552
rect 701 -1576 704 -1574
rect 708 -1576 771 -1574
rect 779 -1576 782 -1574
rect -196 -1580 -193 -1578
rect -189 -1580 -126 -1578
rect -118 -1580 -115 -1578
rect 233 -1579 236 -1577
rect 240 -1579 303 -1577
rect 311 -1579 314 -1577
rect 462 -1579 465 -1577
rect 469 -1579 532 -1577
rect 540 -1579 543 -1577
rect 735 -1631 738 -1629
rect 742 -1631 805 -1629
rect 813 -1631 816 -1629
rect -162 -1635 -159 -1633
rect -155 -1635 -92 -1633
rect -84 -1635 -81 -1633
rect 267 -1634 270 -1632
rect 274 -1634 337 -1632
rect 345 -1634 348 -1632
rect 496 -1634 499 -1632
rect 503 -1634 566 -1632
rect 574 -1634 577 -1632
rect 670 -1638 673 -1636
rect 677 -1638 704 -1636
rect 712 -1638 715 -1636
rect -227 -1642 -224 -1640
rect -220 -1642 -193 -1640
rect -185 -1642 -182 -1640
rect 202 -1641 205 -1639
rect 209 -1641 236 -1639
rect 244 -1641 247 -1639
rect 431 -1641 434 -1639
rect 438 -1641 465 -1639
rect 473 -1641 476 -1639
rect -227 -1667 -224 -1665
rect -220 -1667 -193 -1665
rect -185 -1667 -182 -1665
rect 202 -1666 205 -1664
rect 209 -1666 236 -1664
rect 244 -1666 247 -1664
rect -126 -1671 -123 -1669
rect -119 -1671 -92 -1669
rect -84 -1671 -81 -1669
rect 670 -1663 673 -1661
rect 677 -1663 704 -1661
rect 712 -1663 715 -1661
rect 431 -1666 434 -1664
rect 438 -1666 465 -1664
rect 473 -1666 476 -1664
rect 303 -1670 306 -1668
rect 310 -1670 337 -1668
rect 345 -1670 348 -1668
rect 771 -1667 774 -1665
rect 778 -1667 805 -1665
rect 813 -1667 816 -1665
rect 532 -1670 535 -1668
rect 539 -1670 566 -1668
rect 574 -1670 577 -1668
rect -227 -1692 -224 -1690
rect -220 -1692 -193 -1690
rect -185 -1692 -182 -1690
rect 202 -1691 205 -1689
rect 209 -1691 236 -1689
rect 244 -1691 247 -1689
rect -162 -1696 -159 -1694
rect -155 -1696 -92 -1694
rect -84 -1696 -81 -1694
rect 670 -1688 673 -1686
rect 677 -1688 704 -1686
rect 712 -1688 715 -1686
rect 431 -1691 434 -1689
rect 438 -1691 465 -1689
rect 473 -1691 476 -1689
rect 267 -1695 270 -1693
rect 274 -1695 337 -1693
rect 345 -1695 348 -1693
rect 735 -1692 738 -1690
rect 742 -1692 805 -1690
rect 813 -1692 816 -1690
rect 496 -1695 499 -1693
rect 503 -1695 566 -1693
rect 574 -1695 577 -1693
rect 735 -1717 738 -1715
rect 742 -1717 805 -1715
rect 813 -1717 816 -1715
rect -162 -1721 -159 -1719
rect -155 -1721 -92 -1719
rect -84 -1721 -81 -1719
rect 267 -1720 270 -1718
rect 274 -1720 337 -1718
rect 345 -1720 348 -1718
rect 496 -1720 499 -1718
rect 503 -1720 566 -1718
rect 574 -1720 577 -1718
rect 645 -1733 648 -1731
rect 652 -1733 692 -1731
rect 700 -1733 703 -1731
rect -252 -1737 -249 -1735
rect -245 -1737 -205 -1735
rect -197 -1737 -194 -1735
rect 177 -1736 180 -1734
rect 184 -1736 224 -1734
rect 232 -1736 235 -1734
rect 406 -1736 409 -1734
rect 413 -1736 453 -1734
rect 461 -1736 464 -1734
rect 771 -1742 774 -1740
rect 778 -1742 805 -1740
rect 813 -1742 816 -1740
rect -126 -1746 -123 -1744
rect -119 -1746 -92 -1744
rect -84 -1746 -81 -1744
rect 303 -1745 306 -1743
rect 310 -1745 337 -1743
rect 345 -1745 348 -1743
rect 532 -1745 535 -1743
rect 539 -1745 566 -1743
rect 574 -1745 577 -1743
rect 645 -1758 648 -1756
rect 652 -1758 692 -1756
rect 700 -1758 703 -1756
rect -252 -1762 -249 -1760
rect -245 -1762 -205 -1760
rect -197 -1762 -194 -1760
rect 177 -1761 180 -1759
rect 184 -1761 224 -1759
rect 232 -1761 235 -1759
rect 406 -1761 409 -1759
rect 413 -1761 453 -1759
rect 461 -1761 464 -1759
rect 735 -1767 738 -1765
rect 742 -1767 805 -1765
rect 813 -1767 816 -1765
rect -162 -1771 -159 -1769
rect -155 -1771 -92 -1769
rect -84 -1771 -81 -1769
rect 267 -1770 270 -1768
rect 274 -1770 337 -1768
rect 345 -1770 348 -1768
rect 496 -1770 499 -1768
rect 503 -1770 566 -1768
rect 574 -1770 577 -1768
rect 658 -1783 661 -1781
rect 665 -1783 692 -1781
rect 700 -1783 703 -1781
rect -239 -1787 -236 -1785
rect -232 -1787 -205 -1785
rect -197 -1787 -194 -1785
rect 190 -1786 193 -1784
rect 197 -1786 224 -1784
rect 232 -1786 235 -1784
rect 419 -1786 422 -1784
rect 426 -1786 453 -1784
rect 461 -1786 464 -1784
rect 483 -1911 486 -1909
rect 490 -1911 553 -1909
rect 561 -1911 564 -1909
rect 409 -1918 412 -1916
rect 416 -1918 443 -1916
rect 451 -1918 454 -1916
rect 1 -1922 4 -1920
rect 8 -1922 71 -1920
rect 79 -1922 82 -1920
rect 239 -1922 242 -1920
rect 246 -1922 309 -1920
rect 317 -1922 320 -1920
rect 676 -1919 679 -1917
rect 683 -1919 746 -1917
rect 754 -1919 757 -1917
rect 602 -1926 605 -1924
rect 609 -1926 636 -1924
rect 644 -1926 647 -1924
rect -73 -1929 -70 -1927
rect -66 -1929 -39 -1927
rect -31 -1929 -28 -1927
rect 165 -1929 168 -1927
rect 172 -1929 199 -1927
rect 207 -1929 210 -1927
rect 409 -1943 412 -1941
rect 416 -1943 443 -1941
rect 451 -1943 454 -1941
rect -73 -1954 -70 -1952
rect -66 -1954 -39 -1952
rect -31 -1954 -28 -1952
rect 519 -1947 522 -1945
rect 526 -1947 553 -1945
rect 561 -1947 564 -1945
rect 165 -1954 168 -1952
rect 172 -1954 199 -1952
rect 207 -1954 210 -1952
rect 37 -1958 40 -1956
rect 44 -1958 71 -1956
rect 79 -1958 82 -1956
rect 602 -1951 605 -1949
rect 609 -1951 636 -1949
rect 644 -1951 647 -1949
rect 712 -1955 715 -1953
rect 719 -1955 746 -1953
rect 754 -1955 757 -1953
rect 275 -1958 278 -1956
rect 282 -1958 309 -1956
rect 317 -1958 320 -1956
rect 409 -1968 412 -1966
rect 416 -1968 443 -1966
rect 451 -1968 454 -1966
rect -73 -1979 -70 -1977
rect -66 -1979 -39 -1977
rect -31 -1979 -28 -1977
rect 483 -1972 486 -1970
rect 490 -1972 553 -1970
rect 561 -1972 564 -1970
rect 165 -1979 168 -1977
rect 172 -1979 199 -1977
rect 207 -1979 210 -1977
rect 1 -1983 4 -1981
rect 8 -1983 71 -1981
rect 79 -1983 82 -1981
rect 602 -1976 605 -1974
rect 609 -1976 636 -1974
rect 644 -1976 647 -1974
rect 676 -1980 679 -1978
rect 683 -1980 746 -1978
rect 754 -1980 757 -1978
rect 239 -1983 242 -1981
rect 246 -1983 309 -1981
rect 317 -1983 320 -1981
rect 483 -1997 486 -1995
rect 490 -1997 553 -1995
rect 561 -1997 564 -1995
rect 676 -2005 679 -2003
rect 683 -2005 746 -2003
rect 754 -2005 757 -2003
rect 1 -2008 4 -2006
rect 8 -2008 71 -2006
rect 79 -2008 82 -2006
rect 239 -2008 242 -2006
rect 246 -2008 309 -2006
rect 317 -2008 320 -2006
rect 519 -2022 522 -2020
rect 526 -2022 553 -2020
rect 561 -2022 564 -2020
rect 712 -2030 715 -2028
rect 719 -2030 746 -2028
rect 754 -2030 757 -2028
rect 37 -2033 40 -2031
rect 44 -2033 71 -2031
rect 79 -2033 82 -2031
rect 275 -2033 278 -2031
rect 282 -2033 309 -2031
rect 317 -2033 320 -2031
rect 483 -2047 486 -2045
rect 490 -2047 553 -2045
rect 561 -2047 564 -2045
rect 676 -2055 679 -2053
rect 683 -2055 746 -2053
rect 754 -2055 757 -2053
rect 1 -2058 4 -2056
rect 8 -2058 71 -2056
rect 79 -2058 82 -2056
rect 239 -2058 242 -2056
rect 246 -2058 309 -2056
rect 317 -2058 320 -2056
rect 710 -2110 713 -2108
rect 717 -2110 780 -2108
rect 788 -2110 791 -2108
rect 35 -2113 38 -2111
rect 42 -2113 105 -2111
rect 113 -2113 116 -2111
rect 273 -2113 276 -2111
rect 280 -2113 343 -2111
rect 351 -2113 354 -2111
rect 645 -2117 648 -2115
rect 652 -2117 679 -2115
rect 687 -2117 690 -2115
rect -30 -2120 -27 -2118
rect -23 -2120 4 -2118
rect 12 -2120 15 -2118
rect 208 -2120 211 -2118
rect 215 -2120 242 -2118
rect 250 -2120 253 -2118
rect -30 -2145 -27 -2143
rect -23 -2145 4 -2143
rect 12 -2145 15 -2143
rect 645 -2142 648 -2140
rect 652 -2142 679 -2140
rect 687 -2142 690 -2140
rect 208 -2145 211 -2143
rect 215 -2145 242 -2143
rect 250 -2145 253 -2143
rect 71 -2149 74 -2147
rect 78 -2149 105 -2147
rect 113 -2149 116 -2147
rect 746 -2146 749 -2144
rect 753 -2146 780 -2144
rect 788 -2146 791 -2144
rect 309 -2149 312 -2147
rect 316 -2149 343 -2147
rect 351 -2149 354 -2147
rect -30 -2170 -27 -2168
rect -23 -2170 4 -2168
rect 12 -2170 15 -2168
rect 645 -2167 648 -2165
rect 652 -2167 679 -2165
rect 687 -2167 690 -2165
rect 208 -2170 211 -2168
rect 215 -2170 242 -2168
rect 250 -2170 253 -2168
rect 35 -2174 38 -2172
rect 42 -2174 105 -2172
rect 113 -2174 116 -2172
rect 710 -2171 713 -2169
rect 717 -2171 780 -2169
rect 788 -2171 791 -2169
rect 273 -2174 276 -2172
rect 280 -2174 343 -2172
rect 351 -2174 354 -2172
rect 710 -2196 713 -2194
rect 717 -2196 780 -2194
rect 788 -2196 791 -2194
rect 35 -2199 38 -2197
rect 42 -2199 105 -2197
rect 113 -2199 116 -2197
rect 273 -2199 276 -2197
rect 280 -2199 343 -2197
rect 351 -2199 354 -2197
rect 620 -2212 623 -2210
rect 627 -2212 667 -2210
rect 675 -2212 678 -2210
rect -55 -2215 -52 -2213
rect -48 -2215 -8 -2213
rect 0 -2215 3 -2213
rect 183 -2215 186 -2213
rect 190 -2215 230 -2213
rect 238 -2215 241 -2213
rect 746 -2221 749 -2219
rect 753 -2221 780 -2219
rect 788 -2221 791 -2219
rect 71 -2224 74 -2222
rect 78 -2224 105 -2222
rect 113 -2224 116 -2222
rect 309 -2224 312 -2222
rect 316 -2224 343 -2222
rect 351 -2224 354 -2222
rect 620 -2237 623 -2235
rect 627 -2237 667 -2235
rect 675 -2237 678 -2235
rect -55 -2240 -52 -2238
rect -48 -2240 -8 -2238
rect 0 -2240 3 -2238
rect 183 -2240 186 -2238
rect 190 -2240 230 -2238
rect 238 -2240 241 -2238
rect 710 -2246 713 -2244
rect 717 -2246 780 -2244
rect 788 -2246 791 -2244
rect 35 -2249 38 -2247
rect 42 -2249 105 -2247
rect 113 -2249 116 -2247
rect 273 -2249 276 -2247
rect 280 -2249 343 -2247
rect 351 -2249 354 -2247
rect 633 -2262 636 -2260
rect 640 -2262 667 -2260
rect 675 -2262 678 -2260
rect -42 -2265 -39 -2263
rect -35 -2265 -8 -2263
rect 0 -2265 3 -2263
rect 196 -2265 199 -2263
rect 203 -2265 230 -2263
rect 238 -2265 241 -2263
<< polycontact >>
rect 37 -759 41 -755
rect 97 -759 101 -755
rect 157 -759 161 -755
rect 217 -759 221 -755
rect 277 -759 281 -755
rect 337 -759 341 -755
rect 397 -759 401 -755
rect 457 -759 461 -755
rect 517 -759 521 -755
rect 577 -759 581 -755
rect 637 -759 641 -755
rect 697 -759 701 -755
rect 757 -759 761 -755
rect 817 -759 821 -755
rect 877 -759 881 -755
rect 937 -759 941 -755
rect 28 -784 32 -780
rect 88 -784 92 -780
rect 148 -784 152 -780
rect 208 -784 212 -780
rect 268 -784 272 -780
rect 328 -784 332 -780
rect 388 -784 392 -780
rect 448 -784 452 -780
rect 508 -784 512 -780
rect 568 -784 572 -780
rect 628 -784 632 -780
rect 688 -784 692 -780
rect 748 -784 752 -780
rect 808 -784 812 -780
rect 868 -784 872 -780
rect 928 -784 932 -780
rect 37 -809 41 -805
rect 97 -809 101 -805
rect 157 -809 161 -805
rect 217 -809 221 -805
rect 277 -809 281 -805
rect 337 -809 341 -805
rect 397 -809 401 -805
rect 457 -809 461 -805
rect 517 -809 521 -805
rect 577 -809 581 -805
rect 637 -809 641 -805
rect 697 -809 701 -805
rect 757 -809 761 -805
rect 817 -809 821 -805
rect 877 -809 881 -805
rect 937 -809 941 -805
rect 469 -872 473 -868
rect 359 -879 363 -875
rect 706 -876 710 -872
rect 889 -876 893 -872
rect 596 -883 600 -879
rect 779 -883 783 -879
rect 124 -892 128 -888
rect 14 -899 18 -895
rect 350 -904 354 -900
rect 469 -908 473 -904
rect 587 -908 591 -904
rect 706 -912 710 -908
rect 770 -908 774 -904
rect 889 -912 893 -908
rect 5 -924 9 -920
rect 124 -928 128 -924
rect 359 -929 363 -925
rect 469 -933 473 -929
rect 596 -933 600 -929
rect 706 -937 710 -933
rect 779 -933 783 -929
rect 889 -937 893 -933
rect 14 -949 18 -945
rect 124 -953 128 -949
rect 469 -958 473 -954
rect 706 -962 710 -958
rect 889 -962 893 -958
rect 124 -978 128 -974
rect 469 -983 473 -979
rect 706 -987 710 -983
rect 889 -987 893 -983
rect 124 -1003 128 -999
rect 469 -1008 473 -1004
rect 706 -1012 710 -1008
rect 889 -1012 893 -1008
rect 124 -1028 128 -1024
rect 158 -1083 162 -1079
rect 57 -1090 61 -1086
rect 48 -1115 52 -1111
rect 158 -1119 162 -1115
rect 57 -1140 61 -1136
rect 158 -1144 162 -1140
rect 158 -1169 162 -1165
rect 47 -1185 51 -1181
rect 158 -1194 162 -1190
rect 40 -1210 44 -1206
rect 158 -1219 162 -1215
rect 45 -1235 49 -1231
rect -140 -1442 -136 -1438
rect 289 -1441 293 -1437
rect 518 -1441 522 -1437
rect 757 -1438 761 -1434
rect -250 -1449 -246 -1445
rect 179 -1448 183 -1444
rect 408 -1448 412 -1444
rect 647 -1445 651 -1441
rect -259 -1474 -255 -1470
rect 170 -1473 174 -1469
rect -140 -1478 -136 -1474
rect 289 -1477 293 -1473
rect 399 -1473 403 -1469
rect 638 -1470 642 -1466
rect 518 -1477 522 -1473
rect 757 -1474 761 -1470
rect -250 -1499 -246 -1495
rect 179 -1498 183 -1494
rect -140 -1503 -136 -1499
rect 289 -1502 293 -1498
rect 408 -1498 412 -1494
rect 647 -1495 651 -1491
rect 518 -1502 522 -1498
rect 757 -1499 761 -1495
rect -140 -1528 -136 -1524
rect 289 -1527 293 -1523
rect 518 -1527 522 -1523
rect 757 -1524 761 -1520
rect -140 -1553 -136 -1549
rect 289 -1552 293 -1548
rect 518 -1552 522 -1548
rect 757 -1549 761 -1545
rect -140 -1578 -136 -1574
rect 289 -1577 293 -1573
rect 518 -1577 522 -1573
rect 757 -1574 761 -1570
rect -106 -1633 -102 -1629
rect 323 -1632 327 -1628
rect 552 -1632 556 -1628
rect 791 -1629 795 -1625
rect -207 -1640 -203 -1636
rect 222 -1639 226 -1635
rect 451 -1639 455 -1635
rect 690 -1636 694 -1632
rect -216 -1665 -212 -1661
rect 213 -1664 217 -1660
rect -106 -1669 -102 -1665
rect 323 -1668 327 -1664
rect 442 -1664 446 -1660
rect 681 -1661 685 -1657
rect 552 -1668 556 -1664
rect 791 -1665 795 -1661
rect -207 -1690 -203 -1686
rect 222 -1689 226 -1685
rect -106 -1694 -102 -1690
rect 323 -1693 327 -1689
rect 451 -1689 455 -1685
rect 690 -1686 694 -1682
rect 552 -1693 556 -1689
rect 791 -1690 795 -1686
rect -106 -1719 -102 -1715
rect 323 -1718 327 -1714
rect 552 -1718 556 -1714
rect 791 -1715 795 -1711
rect -217 -1735 -213 -1731
rect 212 -1734 216 -1730
rect 441 -1734 445 -1730
rect 680 -1731 684 -1727
rect -106 -1744 -102 -1740
rect 323 -1743 327 -1739
rect 552 -1743 556 -1739
rect 791 -1740 795 -1736
rect -224 -1760 -220 -1756
rect 205 -1759 209 -1755
rect 434 -1759 438 -1755
rect 673 -1756 677 -1752
rect -106 -1769 -102 -1765
rect 323 -1768 327 -1764
rect 552 -1768 556 -1764
rect 791 -1765 795 -1761
rect -219 -1785 -215 -1781
rect 210 -1784 214 -1780
rect 439 -1784 443 -1780
rect 678 -1781 682 -1777
rect 539 -1909 543 -1905
rect 57 -1920 61 -1916
rect 295 -1920 299 -1916
rect 429 -1916 433 -1912
rect 732 -1917 736 -1913
rect -53 -1927 -49 -1923
rect 185 -1927 189 -1923
rect 622 -1924 626 -1920
rect 420 -1941 424 -1937
rect -62 -1952 -58 -1948
rect 57 -1956 61 -1952
rect 176 -1952 180 -1948
rect 539 -1945 543 -1941
rect 295 -1956 299 -1952
rect 613 -1949 617 -1945
rect 732 -1953 736 -1949
rect 429 -1966 433 -1962
rect -53 -1977 -49 -1973
rect 57 -1981 61 -1977
rect 185 -1977 189 -1973
rect 539 -1970 543 -1966
rect 295 -1981 299 -1977
rect 622 -1974 626 -1970
rect 732 -1978 736 -1974
rect 539 -1995 543 -1991
rect 57 -2006 61 -2002
rect 295 -2006 299 -2002
rect 732 -2003 736 -1999
rect 539 -2020 543 -2016
rect 57 -2031 61 -2027
rect 295 -2031 299 -2027
rect 732 -2028 736 -2024
rect 539 -2045 543 -2041
rect 57 -2056 61 -2052
rect 295 -2056 299 -2052
rect 732 -2053 736 -2049
rect 91 -2111 95 -2107
rect 329 -2111 333 -2107
rect 766 -2108 770 -2104
rect -10 -2118 -6 -2114
rect 228 -2118 232 -2114
rect 665 -2115 669 -2111
rect -19 -2143 -15 -2139
rect 91 -2147 95 -2143
rect 219 -2143 223 -2139
rect 656 -2140 660 -2136
rect 329 -2147 333 -2143
rect 766 -2144 770 -2140
rect -10 -2168 -6 -2164
rect 91 -2172 95 -2168
rect 228 -2168 232 -2164
rect 665 -2165 669 -2161
rect 329 -2172 333 -2168
rect 766 -2169 770 -2165
rect 91 -2197 95 -2193
rect 329 -2197 333 -2193
rect 766 -2194 770 -2190
rect -20 -2213 -16 -2209
rect 218 -2213 222 -2209
rect 655 -2210 659 -2206
rect 91 -2222 95 -2218
rect 329 -2222 333 -2218
rect 766 -2219 770 -2215
rect -27 -2238 -23 -2234
rect 211 -2238 215 -2234
rect 648 -2235 652 -2231
rect 91 -2247 95 -2243
rect 329 -2247 333 -2243
rect 766 -2244 770 -2240
rect -22 -2263 -18 -2259
rect 216 -2263 220 -2259
rect 653 -2260 657 -2256
<< metal1 >>
rect 10 -680 36 -677
rect 41 -680 96 -677
rect 101 -680 276 -677
rect 281 -680 456 -677
rect 10 -688 156 -685
rect 161 -688 336 -685
rect 341 -688 396 -685
rect 401 -688 696 -685
rect 10 -696 216 -693
rect 221 -696 576 -693
rect 581 -696 636 -693
rect 641 -696 816 -693
rect 10 -704 516 -701
rect 521 -704 756 -701
rect 761 -704 876 -701
rect 881 -704 927 -701
rect 10 -714 28 -711
rect 33 -714 147 -711
rect 152 -714 207 -711
rect 212 -714 507 -711
rect 10 -722 87 -719
rect 92 -722 327 -719
rect 332 -722 567 -719
rect 572 -722 747 -719
rect 10 -730 267 -727
rect 272 -730 387 -727
rect 392 -730 627 -727
rect 632 -730 867 -727
rect 10 -738 447 -735
rect 452 -738 687 -735
rect 692 -738 807 -735
rect 812 -738 936 -735
rect 64 -744 999 -741
rect 11 -754 15 -744
rect 11 -758 20 -754
rect 11 -804 15 -758
rect 20 -779 24 -766
rect 28 -780 32 -753
rect 37 -755 41 -752
rect 64 -754 68 -744
rect 59 -758 68 -754
rect 51 -770 59 -766
rect 37 -775 59 -770
rect 37 -787 41 -775
rect 51 -779 59 -775
rect 64 -787 68 -758
rect 24 -791 41 -787
rect 59 -791 68 -787
rect 11 -808 20 -804
rect 37 -805 41 -791
rect 64 -804 68 -791
rect 11 -825 15 -808
rect 59 -808 68 -804
rect 24 -816 51 -812
rect 37 -840 41 -816
rect 64 -823 68 -808
rect 71 -754 75 -748
rect 71 -758 80 -754
rect 71 -804 75 -758
rect 80 -779 84 -766
rect 88 -780 92 -753
rect 97 -755 101 -752
rect 124 -754 128 -744
rect 119 -758 128 -754
rect 111 -770 119 -766
rect 97 -775 119 -770
rect 97 -787 101 -775
rect 111 -779 119 -775
rect 124 -787 128 -758
rect 84 -791 101 -787
rect 119 -791 128 -787
rect 71 -808 80 -804
rect 97 -805 101 -791
rect 124 -804 128 -791
rect 71 -826 75 -808
rect 119 -808 128 -804
rect 84 -816 111 -812
rect -155 -843 41 -840
rect -276 -1444 -272 -1402
rect -155 -1408 -152 -843
rect 97 -859 101 -816
rect 124 -823 128 -808
rect 131 -754 135 -748
rect 131 -758 140 -754
rect 131 -804 135 -758
rect 140 -779 144 -766
rect 148 -780 152 -753
rect 157 -755 161 -752
rect 184 -754 188 -744
rect 179 -758 188 -754
rect 171 -770 179 -766
rect 157 -775 179 -770
rect 157 -787 161 -775
rect 171 -779 179 -775
rect 184 -787 188 -758
rect 144 -791 161 -787
rect 179 -791 188 -787
rect 131 -808 140 -804
rect 157 -805 161 -791
rect 184 -804 188 -791
rect 131 -826 135 -808
rect 179 -808 188 -804
rect 144 -816 171 -812
rect 157 -843 161 -816
rect 184 -823 188 -808
rect 191 -754 195 -748
rect 191 -758 200 -754
rect 191 -804 195 -758
rect 200 -779 204 -766
rect 208 -780 212 -753
rect 217 -755 221 -752
rect 244 -754 248 -744
rect 239 -758 248 -754
rect 231 -770 239 -766
rect 217 -775 239 -770
rect 217 -787 221 -775
rect 231 -779 239 -775
rect 244 -787 248 -758
rect 204 -791 221 -787
rect 239 -791 248 -787
rect 191 -808 200 -804
rect 217 -805 221 -791
rect 244 -804 248 -791
rect 191 -826 195 -808
rect 239 -808 248 -804
rect 204 -816 231 -812
rect 124 -846 161 -843
rect 97 -862 112 -859
rect -12 -894 -8 -867
rect 124 -869 128 -846
rect 5 -872 128 -869
rect -12 -898 -3 -894
rect -12 -944 -8 -898
rect -3 -919 1 -906
rect 5 -920 9 -872
rect 124 -875 128 -872
rect 171 -870 212 -867
rect 124 -878 162 -875
rect 14 -895 18 -880
rect 41 -894 45 -888
rect 36 -898 45 -894
rect 28 -910 36 -906
rect 14 -915 36 -910
rect 14 -927 18 -915
rect 28 -919 36 -915
rect 41 -927 45 -898
rect 1 -931 18 -927
rect 36 -931 45 -927
rect -12 -948 -3 -944
rect 14 -945 18 -931
rect 41 -944 45 -931
rect -12 -1009 -8 -948
rect 36 -948 45 -944
rect 1 -956 13 -952
rect 18 -956 28 -952
rect 41 -958 45 -948
rect 62 -891 71 -887
rect 124 -888 128 -878
rect 151 -887 155 -881
rect 62 -973 65 -891
rect 146 -891 155 -887
rect 75 -899 89 -895
rect 86 -948 89 -899
rect 75 -952 89 -948
rect 75 -960 81 -956
rect 62 -977 71 -973
rect 71 -998 75 -985
rect 71 -1009 75 -1003
rect -12 -1014 75 -1009
rect 31 -1085 35 -1014
rect 71 -1023 75 -1014
rect 78 -1031 81 -960
rect 75 -1035 81 -1031
rect 86 -1045 89 -952
rect 92 -899 138 -895
rect 92 -1031 95 -899
rect 151 -906 155 -896
rect 159 -910 162 -878
rect 124 -913 162 -910
rect 98 -923 102 -917
rect 98 -927 107 -923
rect 124 -924 128 -913
rect 151 -923 155 -922
rect 98 -997 102 -927
rect 146 -927 155 -923
rect 111 -935 138 -931
rect 124 -949 128 -935
rect 151 -948 155 -927
rect 146 -952 155 -948
rect 121 -970 128 -967
rect 118 -992 121 -972
rect 124 -974 128 -970
rect 138 -973 146 -960
rect 151 -967 155 -952
rect 146 -985 161 -981
rect 118 -995 128 -992
rect 103 -1002 107 -998
rect 124 -999 128 -995
rect 150 -998 155 -997
rect 98 -1017 102 -1002
rect 146 -1002 155 -998
rect 111 -1010 138 -1006
rect 124 -1024 128 -1010
rect 151 -1017 155 -1002
rect 158 -1023 161 -985
rect 146 -1027 161 -1023
rect 92 -1035 138 -1031
rect 158 -1045 161 -1027
rect 86 -1048 161 -1045
rect 158 -1066 161 -1048
rect 171 -1058 175 -870
rect 158 -1069 196 -1066
rect 158 -1072 162 -1069
rect 57 -1075 162 -1072
rect 31 -1089 40 -1085
rect 31 -1135 35 -1089
rect 40 -1110 44 -1097
rect 48 -1111 52 -1078
rect 57 -1086 61 -1075
rect 84 -1085 88 -1079
rect 79 -1089 88 -1085
rect 71 -1101 79 -1097
rect 57 -1106 79 -1101
rect 57 -1118 61 -1106
rect 71 -1110 79 -1106
rect 84 -1118 88 -1089
rect 44 -1122 61 -1118
rect 79 -1122 88 -1118
rect 31 -1139 40 -1135
rect 57 -1136 61 -1122
rect 84 -1135 88 -1122
rect 31 -1151 35 -1139
rect 79 -1139 88 -1135
rect 44 -1147 71 -1143
rect 6 -1154 35 -1151
rect 6 -1180 10 -1154
rect 57 -1163 61 -1147
rect 84 -1149 88 -1139
rect 96 -1082 105 -1078
rect 158 -1079 162 -1075
rect 185 -1078 189 -1072
rect 47 -1166 61 -1163
rect 96 -1164 99 -1082
rect 180 -1082 189 -1078
rect 109 -1090 123 -1086
rect 120 -1139 123 -1090
rect 109 -1143 123 -1139
rect 109 -1151 115 -1147
rect 6 -1184 15 -1180
rect 6 -1205 10 -1184
rect 19 -1192 25 -1188
rect 6 -1209 15 -1205
rect 6 -1224 10 -1209
rect 22 -1213 25 -1192
rect 40 -1206 44 -1174
rect 47 -1181 51 -1166
rect 96 -1168 105 -1164
rect 72 -1180 76 -1179
rect 67 -1184 76 -1180
rect 59 -1205 67 -1192
rect 19 -1217 59 -1213
rect 6 -1227 19 -1224
rect 19 -1230 23 -1227
rect 19 -1234 28 -1230
rect 45 -1231 49 -1217
rect 72 -1230 76 -1184
rect 105 -1189 109 -1176
rect 105 -1197 109 -1194
rect 95 -1201 109 -1197
rect 95 -1224 98 -1201
rect 105 -1214 109 -1201
rect 112 -1222 115 -1151
rect 84 -1227 98 -1224
rect 109 -1226 115 -1222
rect 19 -1256 23 -1234
rect 67 -1234 76 -1230
rect 32 -1242 59 -1238
rect 45 -1280 49 -1242
rect 72 -1248 76 -1234
rect 120 -1236 123 -1143
rect 126 -1090 172 -1086
rect 126 -1222 129 -1090
rect 185 -1097 189 -1087
rect 193 -1101 196 -1069
rect 158 -1104 196 -1101
rect 132 -1114 136 -1108
rect 132 -1118 141 -1114
rect 158 -1115 162 -1104
rect 185 -1114 189 -1113
rect 132 -1188 136 -1118
rect 180 -1118 189 -1114
rect 145 -1126 172 -1122
rect 158 -1140 162 -1126
rect 185 -1139 189 -1118
rect 180 -1143 189 -1139
rect 155 -1161 162 -1158
rect 152 -1183 155 -1163
rect 158 -1165 162 -1161
rect 172 -1164 180 -1151
rect 185 -1158 189 -1143
rect 180 -1176 195 -1172
rect 152 -1186 162 -1183
rect 137 -1189 145 -1188
rect 137 -1193 141 -1189
rect 158 -1190 162 -1186
rect 184 -1189 189 -1188
rect 132 -1208 136 -1193
rect 180 -1193 189 -1189
rect 145 -1201 172 -1197
rect 158 -1215 162 -1201
rect 185 -1208 189 -1193
rect 192 -1214 195 -1176
rect 180 -1218 195 -1214
rect 126 -1226 172 -1222
rect 192 -1236 195 -1218
rect 120 -1239 195 -1236
rect 192 -1250 195 -1239
rect -140 -1283 49 -1280
rect 102 -1255 195 -1250
rect -140 -1419 -136 -1283
rect 102 -1301 107 -1255
rect 209 -1260 212 -870
rect 145 -1263 212 -1260
rect -259 -1422 -136 -1419
rect -276 -1448 -267 -1444
rect -276 -1494 -272 -1448
rect -267 -1469 -263 -1456
rect -259 -1470 -255 -1422
rect -140 -1425 -136 -1422
rect 46 -1304 107 -1301
rect -140 -1428 -102 -1425
rect -250 -1445 -246 -1430
rect -223 -1444 -219 -1438
rect -228 -1448 -219 -1444
rect -236 -1460 -228 -1456
rect -250 -1465 -228 -1460
rect -250 -1477 -246 -1465
rect -236 -1469 -228 -1465
rect -223 -1477 -219 -1448
rect -263 -1481 -246 -1477
rect -228 -1481 -219 -1477
rect -276 -1498 -267 -1494
rect -250 -1495 -246 -1481
rect -223 -1494 -219 -1481
rect -276 -1559 -272 -1498
rect -228 -1498 -219 -1494
rect -263 -1506 -251 -1502
rect -246 -1506 -236 -1502
rect -223 -1508 -219 -1498
rect -202 -1441 -193 -1437
rect -140 -1438 -136 -1428
rect -113 -1437 -109 -1431
rect -202 -1523 -199 -1441
rect -118 -1441 -109 -1437
rect -189 -1449 -175 -1445
rect -178 -1498 -175 -1449
rect -189 -1502 -175 -1498
rect -189 -1510 -183 -1506
rect -202 -1527 -193 -1523
rect -193 -1548 -189 -1535
rect -193 -1559 -189 -1553
rect -276 -1564 -189 -1559
rect -233 -1635 -229 -1564
rect -193 -1573 -189 -1564
rect -186 -1581 -183 -1510
rect -189 -1585 -183 -1581
rect -178 -1595 -175 -1502
rect -172 -1449 -126 -1445
rect -172 -1581 -169 -1449
rect -113 -1456 -109 -1446
rect -105 -1460 -102 -1428
rect -140 -1463 -102 -1460
rect -166 -1473 -162 -1467
rect -166 -1477 -157 -1473
rect -140 -1474 -136 -1463
rect -113 -1473 -109 -1472
rect -166 -1547 -162 -1477
rect -118 -1477 -109 -1473
rect -153 -1485 -126 -1481
rect -140 -1499 -136 -1485
rect -113 -1498 -109 -1477
rect -118 -1502 -109 -1498
rect -143 -1520 -136 -1517
rect -146 -1542 -143 -1522
rect -140 -1524 -136 -1520
rect -126 -1523 -118 -1510
rect -113 -1517 -109 -1502
rect -118 -1535 -103 -1531
rect -146 -1545 -136 -1542
rect -161 -1552 -157 -1548
rect -140 -1549 -136 -1545
rect -114 -1548 -109 -1547
rect -166 -1567 -162 -1552
rect -118 -1552 -109 -1548
rect -153 -1560 -126 -1556
rect -140 -1574 -136 -1560
rect -113 -1567 -109 -1552
rect -106 -1573 -103 -1535
rect -118 -1577 -103 -1573
rect -172 -1585 -126 -1581
rect -106 -1595 -103 -1577
rect -178 -1598 -103 -1595
rect -106 -1616 -103 -1598
rect -93 -1597 -55 -1594
rect -93 -1608 -89 -1597
rect -106 -1619 -68 -1616
rect -106 -1622 -102 -1619
rect -207 -1625 -102 -1622
rect -233 -1639 -224 -1635
rect -233 -1685 -229 -1639
rect -224 -1660 -220 -1647
rect -216 -1661 -212 -1628
rect -207 -1636 -203 -1625
rect -180 -1635 -176 -1629
rect -185 -1639 -176 -1635
rect -193 -1651 -185 -1647
rect -207 -1656 -185 -1651
rect -207 -1668 -203 -1656
rect -193 -1660 -185 -1656
rect -180 -1668 -176 -1639
rect -220 -1672 -203 -1668
rect -185 -1672 -176 -1668
rect -233 -1689 -224 -1685
rect -207 -1686 -203 -1672
rect -180 -1685 -176 -1672
rect -233 -1701 -229 -1689
rect -185 -1689 -176 -1685
rect -220 -1697 -193 -1693
rect -258 -1704 -229 -1701
rect -258 -1730 -254 -1704
rect -207 -1713 -203 -1697
rect -180 -1699 -176 -1689
rect -168 -1632 -159 -1628
rect -106 -1629 -102 -1625
rect -79 -1628 -75 -1622
rect -217 -1716 -203 -1713
rect -168 -1714 -165 -1632
rect -84 -1632 -75 -1628
rect -155 -1640 -141 -1636
rect -144 -1689 -141 -1640
rect -155 -1693 -141 -1689
rect -155 -1701 -149 -1697
rect -258 -1734 -249 -1730
rect -258 -1755 -254 -1734
rect -245 -1742 -239 -1738
rect -258 -1759 -249 -1755
rect -258 -1774 -254 -1759
rect -242 -1763 -239 -1742
rect -224 -1756 -220 -1724
rect -217 -1731 -213 -1716
rect -168 -1718 -159 -1714
rect -192 -1730 -188 -1729
rect -197 -1734 -188 -1730
rect -205 -1755 -197 -1742
rect -245 -1767 -205 -1763
rect -258 -1777 -245 -1774
rect -245 -1780 -241 -1777
rect -245 -1784 -236 -1780
rect -219 -1781 -215 -1767
rect -192 -1780 -188 -1734
rect -159 -1739 -155 -1726
rect -159 -1747 -155 -1744
rect -169 -1751 -155 -1747
rect -169 -1774 -166 -1751
rect -159 -1764 -155 -1751
rect -152 -1772 -149 -1701
rect -180 -1777 -166 -1774
rect -155 -1776 -149 -1772
rect -245 -1799 -241 -1784
rect -197 -1784 -188 -1780
rect -232 -1792 -205 -1788
rect -219 -2341 -215 -1792
rect -192 -1799 -188 -1784
rect -144 -1786 -141 -1693
rect -138 -1640 -92 -1636
rect -138 -1772 -135 -1640
rect -79 -1647 -75 -1637
rect -71 -1651 -68 -1619
rect -106 -1654 -68 -1651
rect -132 -1664 -128 -1658
rect -132 -1668 -123 -1664
rect -106 -1665 -102 -1654
rect -79 -1664 -75 -1663
rect -132 -1738 -128 -1668
rect -84 -1668 -75 -1664
rect -119 -1676 -92 -1672
rect -106 -1690 -102 -1676
rect -79 -1689 -75 -1668
rect -84 -1693 -75 -1689
rect -109 -1711 -102 -1708
rect -112 -1733 -109 -1713
rect -106 -1715 -102 -1711
rect -92 -1714 -84 -1701
rect -79 -1708 -75 -1693
rect -84 -1726 -69 -1722
rect -112 -1736 -102 -1733
rect -127 -1739 -119 -1738
rect -127 -1743 -123 -1739
rect -106 -1740 -102 -1736
rect -80 -1739 -75 -1738
rect -132 -1758 -128 -1743
rect -84 -1743 -75 -1739
rect -119 -1751 -92 -1747
rect -106 -1765 -102 -1751
rect -79 -1758 -75 -1743
rect -72 -1764 -69 -1726
rect -84 -1768 -69 -1764
rect -138 -1776 -92 -1772
rect -72 -1786 -69 -1768
rect -144 -1789 -69 -1786
rect -72 -1817 -69 -1789
rect -121 -1820 -69 -1817
rect -121 -2341 -118 -1820
rect -58 -1853 -55 -1597
rect -88 -1856 -55 -1853
rect -88 -2048 -85 -1856
rect -79 -1922 -75 -1880
rect 46 -1883 49 -1304
rect 128 -1858 132 -1280
rect 145 -1812 149 -1263
rect 217 -1276 221 -816
rect 244 -823 248 -808
rect 251 -754 255 -748
rect 251 -758 260 -754
rect 251 -804 255 -758
rect 260 -779 264 -766
rect 268 -780 272 -753
rect 277 -755 281 -752
rect 304 -754 308 -744
rect 299 -758 308 -754
rect 291 -770 299 -766
rect 277 -775 299 -770
rect 277 -787 281 -775
rect 291 -779 299 -775
rect 304 -787 308 -758
rect 264 -791 281 -787
rect 299 -791 308 -787
rect 251 -808 260 -804
rect 277 -805 281 -791
rect 304 -804 308 -791
rect 251 -826 255 -808
rect 299 -808 308 -804
rect 264 -816 291 -812
rect 277 -849 281 -816
rect 304 -823 308 -808
rect 311 -754 315 -748
rect 311 -758 320 -754
rect 311 -804 315 -758
rect 320 -779 324 -766
rect 328 -780 332 -753
rect 337 -755 341 -752
rect 364 -754 368 -744
rect 359 -758 368 -754
rect 351 -770 359 -766
rect 337 -775 359 -770
rect 337 -787 341 -775
rect 351 -779 359 -775
rect 364 -787 368 -758
rect 324 -791 341 -787
rect 359 -791 368 -787
rect 311 -808 320 -804
rect 337 -805 341 -791
rect 364 -804 368 -791
rect 311 -826 315 -808
rect 359 -808 368 -804
rect 324 -816 351 -812
rect 337 -848 341 -816
rect 364 -823 368 -808
rect 371 -754 375 -748
rect 371 -758 380 -754
rect 371 -804 375 -758
rect 380 -779 384 -766
rect 388 -780 392 -753
rect 397 -755 401 -752
rect 424 -754 428 -744
rect 419 -758 428 -754
rect 411 -770 419 -766
rect 397 -775 419 -770
rect 397 -787 401 -775
rect 411 -779 419 -775
rect 424 -787 428 -758
rect 384 -791 401 -787
rect 419 -791 428 -787
rect 371 -808 380 -804
rect 397 -805 401 -791
rect 424 -804 428 -791
rect 371 -826 375 -808
rect 419 -808 428 -804
rect 384 -816 411 -812
rect 397 -835 401 -816
rect 424 -823 428 -808
rect 431 -754 435 -748
rect 431 -758 440 -754
rect 431 -804 435 -758
rect 440 -779 444 -766
rect 448 -780 452 -753
rect 457 -755 461 -752
rect 484 -754 488 -744
rect 479 -758 488 -754
rect 471 -770 479 -766
rect 457 -775 479 -770
rect 457 -787 461 -775
rect 471 -779 479 -775
rect 484 -787 488 -758
rect 444 -791 461 -787
rect 479 -791 488 -787
rect 431 -808 440 -804
rect 457 -805 461 -791
rect 484 -804 488 -791
rect 431 -826 435 -808
rect 479 -808 488 -804
rect 444 -816 471 -812
rect 457 -840 461 -816
rect 484 -823 488 -808
rect 491 -754 495 -748
rect 491 -758 500 -754
rect 491 -804 495 -758
rect 500 -779 504 -766
rect 508 -780 512 -753
rect 517 -755 521 -752
rect 544 -754 548 -744
rect 539 -758 548 -754
rect 531 -770 539 -766
rect 517 -775 539 -770
rect 517 -787 521 -775
rect 531 -779 539 -775
rect 544 -787 548 -758
rect 504 -791 521 -787
rect 539 -791 548 -787
rect 491 -808 500 -804
rect 517 -805 521 -791
rect 544 -804 548 -791
rect 491 -826 495 -808
rect 539 -808 548 -804
rect 504 -816 531 -812
rect 517 -839 521 -816
rect 544 -823 548 -808
rect 551 -754 555 -748
rect 551 -758 560 -754
rect 551 -804 555 -758
rect 560 -779 564 -766
rect 568 -780 572 -753
rect 577 -755 581 -752
rect 604 -754 608 -744
rect 599 -758 608 -754
rect 591 -770 599 -766
rect 577 -775 599 -770
rect 577 -787 581 -775
rect 591 -779 599 -775
rect 604 -787 608 -758
rect 564 -791 581 -787
rect 599 -791 608 -787
rect 551 -808 560 -804
rect 577 -805 581 -791
rect 604 -804 608 -791
rect 551 -826 555 -808
rect 599 -808 608 -804
rect 564 -816 591 -812
rect 577 -835 581 -816
rect 604 -823 608 -808
rect 611 -754 615 -748
rect 611 -758 620 -754
rect 611 -804 615 -758
rect 620 -779 624 -766
rect 628 -780 632 -753
rect 637 -755 641 -752
rect 664 -754 668 -744
rect 659 -758 668 -754
rect 651 -770 659 -766
rect 637 -775 659 -770
rect 637 -787 641 -775
rect 651 -779 659 -775
rect 664 -787 668 -758
rect 624 -791 641 -787
rect 659 -791 668 -787
rect 611 -808 620 -804
rect 637 -805 641 -791
rect 664 -804 668 -791
rect 611 -826 615 -808
rect 659 -808 668 -804
rect 624 -816 651 -812
rect 637 -832 641 -816
rect 664 -823 668 -808
rect 671 -754 675 -748
rect 671 -758 680 -754
rect 671 -804 675 -758
rect 680 -779 684 -766
rect 688 -780 692 -753
rect 697 -755 701 -752
rect 724 -754 728 -744
rect 719 -758 728 -754
rect 711 -770 719 -766
rect 697 -775 719 -770
rect 697 -787 701 -775
rect 711 -779 719 -775
rect 724 -787 728 -758
rect 684 -791 701 -787
rect 719 -791 728 -787
rect 671 -808 680 -804
rect 697 -805 701 -791
rect 724 -804 728 -791
rect 671 -826 675 -808
rect 719 -808 728 -804
rect 684 -816 711 -812
rect 697 -832 701 -816
rect 724 -823 728 -808
rect 731 -754 735 -748
rect 731 -758 740 -754
rect 731 -804 735 -758
rect 740 -779 744 -766
rect 748 -780 752 -753
rect 757 -755 761 -752
rect 784 -754 788 -744
rect 779 -758 788 -754
rect 771 -770 779 -766
rect 757 -775 779 -770
rect 757 -787 761 -775
rect 771 -779 779 -775
rect 784 -787 788 -758
rect 744 -791 761 -787
rect 779 -791 788 -787
rect 731 -808 740 -804
rect 757 -805 761 -791
rect 784 -804 788 -791
rect 731 -826 735 -808
rect 779 -808 788 -804
rect 744 -816 771 -812
rect 457 -843 473 -840
rect 517 -842 529 -839
rect 274 -852 281 -849
rect 289 -851 341 -848
rect 469 -849 473 -843
rect 557 -839 581 -835
rect 634 -836 641 -832
rect 694 -836 701 -832
rect 757 -835 761 -816
rect 784 -823 788 -808
rect 791 -754 795 -748
rect 791 -758 800 -754
rect 791 -804 795 -758
rect 800 -779 804 -766
rect 808 -780 812 -753
rect 817 -755 821 -752
rect 844 -754 848 -744
rect 839 -758 848 -754
rect 831 -770 839 -766
rect 817 -775 839 -770
rect 817 -787 821 -775
rect 831 -779 839 -775
rect 844 -787 848 -758
rect 804 -791 821 -787
rect 839 -791 848 -787
rect 791 -808 800 -804
rect 817 -805 821 -791
rect 844 -804 848 -791
rect 791 -826 795 -808
rect 839 -808 848 -804
rect 804 -816 831 -812
rect 634 -839 638 -836
rect 694 -844 698 -836
rect 753 -838 761 -835
rect 694 -847 710 -844
rect 753 -847 757 -838
rect 817 -840 821 -816
rect 844 -823 848 -808
rect 851 -754 855 -748
rect 851 -758 860 -754
rect 851 -804 855 -758
rect 860 -779 864 -766
rect 868 -780 872 -753
rect 877 -755 881 -752
rect 904 -754 908 -744
rect 964 -745 999 -744
rect 899 -758 908 -754
rect 891 -770 899 -766
rect 877 -775 899 -770
rect 877 -787 881 -775
rect 891 -779 899 -775
rect 904 -787 908 -758
rect 864 -791 881 -787
rect 899 -791 908 -787
rect 851 -808 860 -804
rect 877 -805 881 -791
rect 904 -804 908 -791
rect 851 -826 855 -808
rect 899 -808 908 -804
rect 864 -816 891 -812
rect 877 -845 881 -816
rect 904 -823 908 -808
rect 911 -754 915 -748
rect 911 -758 920 -754
rect 911 -804 915 -758
rect 920 -779 924 -766
rect 928 -780 932 -753
rect 937 -755 941 -752
rect 964 -754 968 -745
rect 959 -758 968 -754
rect 951 -770 959 -766
rect 937 -775 959 -770
rect 937 -787 941 -775
rect 951 -779 959 -775
rect 964 -787 968 -758
rect 924 -791 941 -787
rect 959 -791 968 -787
rect 911 -808 920 -804
rect 937 -805 941 -791
rect 964 -804 968 -791
rect 911 -826 915 -808
rect 959 -808 968 -804
rect 924 -816 951 -812
rect 153 -1443 157 -1401
rect 274 -1407 277 -852
rect 289 -1418 293 -851
rect 350 -852 473 -849
rect 333 -874 337 -868
rect 333 -878 342 -874
rect 333 -924 337 -878
rect 342 -899 346 -886
rect 350 -900 354 -852
rect 469 -855 473 -852
rect 706 -853 710 -847
rect 469 -858 507 -855
rect 359 -875 363 -860
rect 386 -874 390 -868
rect 381 -878 390 -874
rect 373 -890 381 -886
rect 359 -895 381 -890
rect 359 -907 363 -895
rect 373 -899 381 -895
rect 386 -907 390 -878
rect 346 -911 363 -907
rect 381 -911 390 -907
rect 333 -928 342 -924
rect 359 -925 363 -911
rect 386 -924 390 -911
rect 333 -970 337 -928
rect 381 -928 390 -924
rect 346 -936 358 -932
rect 363 -936 373 -932
rect 386 -938 390 -928
rect 407 -871 416 -867
rect 469 -868 473 -858
rect 496 -867 500 -861
rect 407 -953 410 -871
rect 491 -871 500 -867
rect 420 -879 434 -875
rect 431 -928 434 -879
rect 420 -932 434 -928
rect 420 -940 426 -936
rect 407 -957 416 -953
rect 416 -970 420 -965
rect 333 -975 373 -970
rect 379 -975 420 -970
rect 416 -978 420 -975
rect 170 -1421 293 -1418
rect 153 -1447 162 -1443
rect 153 -1493 157 -1447
rect 162 -1468 166 -1455
rect 170 -1469 174 -1421
rect 289 -1424 293 -1421
rect 289 -1427 327 -1424
rect 179 -1444 183 -1429
rect 206 -1443 210 -1437
rect 201 -1447 210 -1443
rect 193 -1459 201 -1455
rect 179 -1464 201 -1459
rect 179 -1476 183 -1464
rect 193 -1468 201 -1464
rect 206 -1476 210 -1447
rect 166 -1480 183 -1476
rect 201 -1480 210 -1476
rect 153 -1497 162 -1493
rect 179 -1494 183 -1480
rect 206 -1493 210 -1480
rect 153 -1558 157 -1497
rect 201 -1497 210 -1493
rect 166 -1505 178 -1501
rect 183 -1505 193 -1501
rect 206 -1507 210 -1497
rect 227 -1440 236 -1436
rect 289 -1437 293 -1427
rect 316 -1436 320 -1430
rect 227 -1522 230 -1440
rect 311 -1440 320 -1436
rect 240 -1448 254 -1444
rect 251 -1497 254 -1448
rect 240 -1501 254 -1497
rect 240 -1509 246 -1505
rect 227 -1526 236 -1522
rect 236 -1547 240 -1534
rect 236 -1558 240 -1552
rect 153 -1563 240 -1558
rect 196 -1634 200 -1563
rect 236 -1572 240 -1563
rect 243 -1580 246 -1509
rect 240 -1584 246 -1580
rect 251 -1594 254 -1501
rect 257 -1448 303 -1444
rect 257 -1580 260 -1448
rect 316 -1455 320 -1445
rect 324 -1459 327 -1427
rect 289 -1462 327 -1459
rect 263 -1472 267 -1466
rect 263 -1476 272 -1472
rect 289 -1473 293 -1462
rect 316 -1472 320 -1471
rect 263 -1546 267 -1476
rect 311 -1476 320 -1472
rect 276 -1484 303 -1480
rect 289 -1498 293 -1484
rect 316 -1497 320 -1476
rect 311 -1501 320 -1497
rect 286 -1519 293 -1516
rect 283 -1541 286 -1521
rect 289 -1523 293 -1519
rect 303 -1522 311 -1509
rect 316 -1516 320 -1501
rect 311 -1534 326 -1530
rect 283 -1544 293 -1541
rect 268 -1551 272 -1547
rect 289 -1548 293 -1544
rect 315 -1547 320 -1546
rect 263 -1566 267 -1551
rect 311 -1551 320 -1547
rect 276 -1559 303 -1555
rect 289 -1573 293 -1559
rect 316 -1566 320 -1551
rect 323 -1572 326 -1534
rect 311 -1576 326 -1572
rect 257 -1584 303 -1580
rect 323 -1594 326 -1576
rect 251 -1597 326 -1594
rect 323 -1615 326 -1597
rect 336 -1607 340 -991
rect 416 -1003 420 -983
rect 423 -1011 426 -940
rect 420 -1015 426 -1011
rect 431 -1025 434 -932
rect 437 -879 483 -875
rect 437 -1011 440 -879
rect 496 -886 500 -876
rect 504 -890 507 -858
rect 587 -856 710 -853
rect 877 -848 893 -845
rect 889 -853 893 -848
rect 469 -893 507 -890
rect 570 -878 574 -872
rect 570 -882 579 -878
rect 443 -903 447 -897
rect 443 -907 452 -903
rect 469 -904 473 -893
rect 496 -903 500 -902
rect 443 -977 447 -907
rect 491 -907 500 -903
rect 456 -915 483 -911
rect 469 -929 473 -915
rect 496 -928 500 -907
rect 491 -932 500 -928
rect 466 -950 473 -947
rect 463 -972 466 -952
rect 469 -954 473 -950
rect 483 -953 491 -940
rect 496 -947 500 -932
rect 570 -928 574 -882
rect 579 -903 583 -890
rect 587 -904 591 -856
rect 706 -859 710 -856
rect 770 -856 893 -853
rect 706 -862 744 -859
rect 596 -879 600 -864
rect 623 -878 627 -872
rect 618 -882 627 -878
rect 610 -894 618 -890
rect 596 -899 618 -894
rect 596 -911 600 -899
rect 610 -903 618 -899
rect 623 -911 627 -882
rect 583 -915 600 -911
rect 618 -915 627 -911
rect 570 -932 579 -928
rect 596 -929 600 -915
rect 623 -928 627 -915
rect 491 -965 506 -961
rect 463 -975 473 -972
rect 448 -982 452 -978
rect 469 -979 473 -975
rect 495 -978 500 -977
rect 443 -997 447 -982
rect 491 -982 500 -978
rect 456 -990 483 -986
rect 469 -1004 473 -990
rect 496 -997 500 -982
rect 503 -1003 506 -965
rect 570 -974 574 -932
rect 618 -932 627 -928
rect 583 -940 595 -936
rect 600 -940 610 -936
rect 623 -942 627 -932
rect 644 -875 653 -871
rect 706 -872 710 -862
rect 733 -871 737 -865
rect 644 -957 647 -875
rect 728 -875 737 -871
rect 657 -883 671 -879
rect 668 -932 671 -883
rect 657 -936 671 -932
rect 657 -944 663 -940
rect 644 -961 653 -957
rect 653 -974 657 -969
rect 570 -979 607 -974
rect 612 -979 657 -974
rect 653 -982 657 -979
rect 491 -1007 506 -1003
rect 437 -1015 483 -1011
rect 503 -1025 506 -1007
rect 653 -1007 657 -987
rect 660 -1015 663 -944
rect 657 -1019 663 -1015
rect 431 -1028 506 -1025
rect 366 -1034 396 -1031
rect 382 -1443 386 -1401
rect 503 -1407 506 -1028
rect 668 -1029 671 -936
rect 674 -883 720 -879
rect 674 -1015 677 -883
rect 733 -890 737 -880
rect 741 -894 744 -862
rect 706 -897 744 -894
rect 753 -878 757 -872
rect 753 -882 762 -878
rect 680 -907 684 -901
rect 680 -911 689 -907
rect 706 -908 710 -897
rect 733 -907 737 -906
rect 680 -981 684 -911
rect 728 -911 737 -907
rect 693 -919 720 -915
rect 706 -933 710 -919
rect 733 -932 737 -911
rect 728 -936 737 -932
rect 703 -954 710 -951
rect 700 -976 703 -956
rect 706 -958 710 -954
rect 720 -957 728 -944
rect 733 -951 737 -936
rect 753 -928 757 -882
rect 762 -903 766 -890
rect 770 -904 774 -856
rect 889 -859 893 -856
rect 889 -862 927 -859
rect 779 -879 783 -864
rect 806 -878 810 -872
rect 801 -882 810 -878
rect 793 -894 801 -890
rect 779 -899 801 -894
rect 779 -911 783 -899
rect 793 -903 801 -899
rect 806 -911 810 -882
rect 766 -915 783 -911
rect 801 -915 810 -911
rect 753 -932 762 -928
rect 779 -929 783 -915
rect 806 -928 810 -915
rect 728 -969 743 -965
rect 700 -979 710 -976
rect 685 -986 689 -982
rect 706 -983 710 -979
rect 732 -982 737 -981
rect 680 -1001 684 -986
rect 728 -986 737 -982
rect 693 -994 720 -990
rect 706 -1008 710 -994
rect 733 -1001 737 -986
rect 740 -1007 743 -969
rect 753 -974 757 -932
rect 801 -932 810 -928
rect 766 -940 778 -936
rect 783 -940 793 -936
rect 806 -942 810 -932
rect 827 -875 836 -871
rect 889 -872 893 -862
rect 916 -871 920 -865
rect 827 -957 830 -875
rect 911 -875 920 -871
rect 840 -883 854 -879
rect 851 -932 854 -883
rect 840 -936 854 -932
rect 840 -944 846 -940
rect 827 -961 836 -957
rect 836 -974 840 -969
rect 753 -979 794 -974
rect 799 -979 840 -974
rect 836 -982 840 -979
rect 728 -1011 743 -1007
rect 836 -1007 840 -987
rect 674 -1019 720 -1015
rect 740 -1029 743 -1011
rect 843 -1015 846 -944
rect 840 -1019 846 -1015
rect 516 -1038 632 -1031
rect 668 -1032 743 -1029
rect 851 -1029 854 -936
rect 857 -883 903 -879
rect 857 -1015 860 -883
rect 916 -890 920 -880
rect 924 -894 927 -862
rect 889 -897 927 -894
rect 863 -907 867 -901
rect 863 -911 872 -907
rect 889 -908 893 -897
rect 916 -907 920 -906
rect 863 -981 867 -911
rect 911 -911 920 -907
rect 876 -919 903 -915
rect 889 -933 893 -919
rect 916 -932 920 -911
rect 911 -936 920 -932
rect 886 -954 893 -951
rect 883 -976 886 -956
rect 889 -958 893 -954
rect 903 -957 911 -944
rect 916 -951 920 -936
rect 911 -969 926 -965
rect 883 -979 893 -976
rect 868 -986 872 -982
rect 889 -983 893 -979
rect 915 -982 920 -981
rect 863 -1001 867 -986
rect 911 -986 920 -982
rect 876 -994 903 -990
rect 889 -1008 893 -994
rect 916 -1001 920 -986
rect 923 -1007 926 -969
rect 911 -1011 926 -1007
rect 857 -1019 903 -1015
rect 923 -1029 926 -1011
rect 851 -1032 926 -1029
rect 535 -1365 608 -1362
rect 399 -1421 516 -1418
rect 382 -1447 391 -1443
rect 382 -1493 386 -1447
rect 391 -1468 395 -1455
rect 399 -1469 403 -1421
rect 518 -1424 522 -1421
rect 408 -1444 412 -1429
rect 518 -1427 556 -1424
rect 435 -1443 439 -1437
rect 430 -1447 439 -1443
rect 422 -1459 430 -1455
rect 408 -1464 430 -1459
rect 408 -1476 412 -1464
rect 422 -1468 430 -1464
rect 435 -1476 439 -1447
rect 395 -1480 412 -1476
rect 430 -1480 439 -1476
rect 382 -1497 391 -1493
rect 408 -1494 412 -1480
rect 435 -1493 439 -1480
rect 382 -1558 386 -1497
rect 430 -1497 439 -1493
rect 395 -1505 407 -1501
rect 412 -1505 422 -1501
rect 435 -1507 439 -1497
rect 456 -1440 465 -1436
rect 518 -1437 522 -1427
rect 545 -1436 549 -1430
rect 456 -1522 459 -1440
rect 540 -1440 549 -1436
rect 469 -1448 483 -1444
rect 480 -1497 483 -1448
rect 469 -1501 483 -1497
rect 469 -1509 475 -1505
rect 456 -1526 465 -1522
rect 465 -1547 469 -1534
rect 465 -1558 469 -1552
rect 382 -1563 469 -1558
rect 323 -1618 361 -1615
rect 323 -1621 327 -1618
rect 222 -1624 327 -1621
rect 196 -1638 205 -1634
rect 196 -1684 200 -1638
rect 205 -1659 209 -1646
rect 213 -1660 217 -1627
rect 222 -1635 226 -1624
rect 249 -1634 253 -1628
rect 244 -1638 253 -1634
rect 236 -1650 244 -1646
rect 222 -1655 244 -1650
rect 222 -1667 226 -1655
rect 236 -1659 244 -1655
rect 249 -1667 253 -1638
rect 209 -1671 226 -1667
rect 244 -1671 253 -1667
rect 196 -1688 205 -1684
rect 222 -1685 226 -1671
rect 249 -1684 253 -1671
rect 196 -1700 200 -1688
rect 244 -1688 253 -1684
rect 209 -1696 236 -1692
rect 171 -1703 200 -1700
rect 171 -1729 175 -1703
rect 222 -1712 226 -1696
rect 249 -1698 253 -1688
rect 261 -1631 270 -1627
rect 323 -1628 327 -1624
rect 350 -1627 354 -1621
rect 212 -1715 226 -1712
rect 261 -1713 264 -1631
rect 345 -1631 354 -1627
rect 274 -1639 288 -1635
rect 285 -1688 288 -1639
rect 274 -1692 288 -1688
rect 274 -1700 280 -1696
rect 171 -1733 180 -1729
rect 171 -1754 175 -1733
rect 184 -1741 190 -1737
rect 171 -1758 180 -1754
rect 171 -1773 175 -1758
rect 187 -1762 190 -1741
rect 205 -1755 209 -1723
rect 212 -1730 216 -1715
rect 261 -1717 270 -1713
rect 237 -1729 241 -1728
rect 232 -1733 241 -1729
rect 224 -1754 232 -1741
rect 184 -1766 224 -1762
rect 171 -1776 184 -1773
rect 184 -1779 188 -1776
rect 184 -1783 193 -1779
rect 210 -1780 214 -1766
rect 237 -1779 241 -1733
rect 270 -1738 274 -1725
rect 270 -1746 274 -1743
rect 260 -1750 274 -1746
rect 260 -1773 263 -1750
rect 270 -1763 274 -1750
rect 277 -1771 280 -1700
rect 249 -1776 263 -1773
rect 274 -1775 280 -1771
rect 184 -1798 188 -1783
rect 232 -1783 241 -1779
rect 197 -1791 224 -1787
rect 210 -1812 214 -1791
rect 237 -1798 241 -1783
rect 285 -1785 288 -1692
rect 291 -1639 337 -1635
rect 291 -1771 294 -1639
rect 350 -1646 354 -1636
rect 358 -1650 361 -1618
rect 323 -1653 361 -1650
rect 425 -1634 429 -1563
rect 465 -1572 469 -1563
rect 472 -1580 475 -1509
rect 469 -1584 475 -1580
rect 480 -1594 483 -1501
rect 486 -1448 532 -1444
rect 486 -1580 489 -1448
rect 545 -1455 549 -1445
rect 553 -1459 556 -1427
rect 518 -1462 556 -1459
rect 492 -1472 496 -1466
rect 492 -1476 501 -1472
rect 518 -1473 522 -1462
rect 545 -1472 549 -1471
rect 492 -1546 496 -1476
rect 540 -1476 549 -1472
rect 505 -1484 532 -1480
rect 518 -1498 522 -1484
rect 545 -1497 549 -1476
rect 540 -1501 549 -1497
rect 515 -1519 522 -1516
rect 512 -1541 515 -1521
rect 518 -1523 522 -1519
rect 532 -1522 540 -1509
rect 545 -1516 549 -1501
rect 540 -1534 555 -1530
rect 512 -1544 522 -1541
rect 497 -1551 501 -1547
rect 518 -1548 522 -1544
rect 544 -1547 549 -1546
rect 492 -1566 496 -1551
rect 540 -1551 549 -1547
rect 505 -1559 532 -1555
rect 518 -1573 522 -1559
rect 545 -1566 549 -1551
rect 552 -1572 555 -1534
rect 540 -1576 555 -1572
rect 486 -1584 532 -1580
rect 552 -1594 555 -1576
rect 480 -1597 555 -1594
rect 552 -1615 555 -1597
rect 565 -1607 569 -1422
rect 552 -1618 590 -1615
rect 552 -1621 556 -1618
rect 451 -1624 556 -1621
rect 425 -1638 434 -1634
rect 297 -1663 301 -1657
rect 297 -1667 306 -1663
rect 323 -1664 327 -1653
rect 350 -1663 354 -1662
rect 297 -1737 301 -1667
rect 345 -1667 354 -1663
rect 310 -1675 337 -1671
rect 323 -1689 327 -1675
rect 350 -1688 354 -1667
rect 345 -1692 354 -1688
rect 320 -1710 327 -1707
rect 317 -1732 320 -1712
rect 323 -1714 327 -1710
rect 337 -1713 345 -1700
rect 350 -1707 354 -1692
rect 425 -1684 429 -1638
rect 434 -1659 438 -1646
rect 442 -1660 446 -1627
rect 451 -1635 455 -1624
rect 478 -1634 482 -1628
rect 473 -1638 482 -1634
rect 465 -1650 473 -1646
rect 451 -1655 473 -1650
rect 451 -1667 455 -1655
rect 465 -1659 473 -1655
rect 478 -1667 482 -1638
rect 438 -1671 455 -1667
rect 473 -1671 482 -1667
rect 425 -1688 434 -1684
rect 451 -1685 455 -1671
rect 478 -1684 482 -1671
rect 425 -1700 429 -1688
rect 473 -1688 482 -1684
rect 438 -1696 465 -1692
rect 400 -1703 429 -1700
rect 345 -1725 360 -1721
rect 317 -1735 327 -1732
rect 302 -1738 310 -1737
rect 302 -1742 306 -1738
rect 323 -1739 327 -1735
rect 349 -1738 354 -1737
rect 297 -1757 301 -1742
rect 345 -1742 354 -1738
rect 310 -1750 337 -1746
rect 323 -1764 327 -1750
rect 350 -1757 354 -1742
rect 357 -1763 360 -1725
rect 345 -1767 360 -1763
rect 291 -1775 337 -1771
rect 357 -1785 360 -1767
rect 400 -1729 404 -1703
rect 451 -1712 455 -1696
rect 478 -1698 482 -1688
rect 490 -1631 499 -1627
rect 552 -1628 556 -1624
rect 579 -1627 583 -1621
rect 441 -1715 455 -1712
rect 490 -1713 493 -1631
rect 574 -1631 583 -1627
rect 503 -1639 517 -1635
rect 514 -1688 517 -1639
rect 503 -1692 517 -1688
rect 503 -1700 509 -1696
rect 400 -1733 409 -1729
rect 400 -1754 404 -1733
rect 413 -1741 419 -1737
rect 400 -1758 409 -1754
rect 400 -1773 404 -1758
rect 416 -1762 419 -1741
rect 434 -1755 438 -1723
rect 441 -1730 445 -1715
rect 490 -1717 499 -1713
rect 466 -1729 470 -1728
rect 461 -1733 470 -1729
rect 453 -1754 461 -1741
rect 413 -1766 453 -1762
rect 400 -1776 413 -1773
rect 285 -1788 360 -1785
rect 145 -1815 214 -1812
rect 357 -1818 360 -1788
rect 413 -1779 417 -1776
rect 413 -1783 422 -1779
rect 439 -1780 443 -1766
rect 466 -1779 470 -1733
rect 499 -1738 503 -1725
rect 499 -1746 503 -1743
rect 489 -1750 503 -1746
rect 489 -1773 492 -1750
rect 499 -1763 503 -1750
rect 506 -1771 509 -1700
rect 478 -1776 492 -1773
rect 503 -1775 509 -1771
rect 413 -1798 417 -1783
rect 461 -1783 470 -1779
rect 426 -1791 453 -1787
rect 330 -1821 360 -1818
rect 128 -1862 287 -1858
rect -62 -1900 61 -1897
rect -79 -1926 -70 -1922
rect -79 -1972 -75 -1926
rect -70 -1947 -66 -1934
rect -62 -1948 -58 -1900
rect 57 -1903 61 -1900
rect 57 -1906 152 -1903
rect -53 -1923 -49 -1908
rect -26 -1922 -22 -1916
rect -31 -1926 -22 -1922
rect -39 -1938 -31 -1934
rect -53 -1943 -31 -1938
rect -53 -1955 -49 -1943
rect -39 -1947 -31 -1943
rect -26 -1955 -22 -1926
rect -66 -1959 -49 -1955
rect -31 -1959 -22 -1955
rect -79 -1976 -70 -1972
rect -53 -1973 -49 -1959
rect -26 -1972 -22 -1959
rect -79 -2037 -75 -1976
rect -31 -1976 -22 -1972
rect -66 -1984 -54 -1980
rect -49 -1984 -39 -1980
rect -26 -1986 -22 -1976
rect -5 -1919 4 -1915
rect 57 -1916 61 -1906
rect 84 -1915 88 -1909
rect -5 -2001 -2 -1919
rect 79 -1919 88 -1915
rect 8 -1927 22 -1923
rect 19 -1976 22 -1927
rect 8 -1980 22 -1976
rect 8 -1988 14 -1984
rect -5 -2005 4 -2001
rect 4 -2026 8 -2013
rect 4 -2037 8 -2031
rect -79 -2042 8 -2037
rect -88 -2052 -70 -2048
rect -73 -2278 -70 -2052
rect -36 -2113 -32 -2042
rect 4 -2051 8 -2042
rect 11 -2059 14 -1988
rect 8 -2063 14 -2059
rect 19 -2073 22 -1980
rect 25 -1927 71 -1923
rect 25 -2059 28 -1927
rect 84 -1934 88 -1924
rect 92 -1938 95 -1906
rect 57 -1941 95 -1938
rect 31 -1951 35 -1945
rect 31 -1955 40 -1951
rect 57 -1952 61 -1941
rect 84 -1951 88 -1950
rect 31 -2025 35 -1955
rect 79 -1955 88 -1951
rect 44 -1963 71 -1959
rect 57 -1977 61 -1963
rect 84 -1976 88 -1955
rect 79 -1980 88 -1976
rect 54 -1998 61 -1995
rect 51 -2020 54 -2000
rect 57 -2002 61 -1998
rect 71 -2001 79 -1988
rect 84 -1995 88 -1980
rect 79 -2013 94 -2009
rect 51 -2023 61 -2020
rect 36 -2030 40 -2026
rect 57 -2027 61 -2023
rect 83 -2026 88 -2025
rect 31 -2045 35 -2030
rect 79 -2030 88 -2026
rect 44 -2038 71 -2034
rect 57 -2052 61 -2038
rect 84 -2045 88 -2030
rect 91 -2051 94 -2013
rect 79 -2055 94 -2051
rect 25 -2063 71 -2059
rect 91 -2073 94 -2055
rect 19 -2076 94 -2073
rect 91 -2094 94 -2076
rect 104 -2073 141 -2070
rect 104 -2086 108 -2073
rect 91 -2097 129 -2094
rect 91 -2100 95 -2097
rect -10 -2103 95 -2100
rect -36 -2117 -27 -2113
rect -36 -2163 -32 -2117
rect -27 -2138 -23 -2125
rect -19 -2139 -15 -2106
rect -10 -2114 -6 -2103
rect 17 -2113 21 -2107
rect 12 -2117 21 -2113
rect 4 -2129 12 -2125
rect -10 -2134 12 -2129
rect -10 -2146 -6 -2134
rect 4 -2138 12 -2134
rect 17 -2146 21 -2117
rect -23 -2150 -6 -2146
rect 12 -2150 21 -2146
rect -36 -2167 -27 -2163
rect -10 -2164 -6 -2150
rect 17 -2163 21 -2150
rect -36 -2179 -32 -2167
rect 12 -2167 21 -2163
rect -23 -2175 4 -2171
rect -61 -2182 -32 -2179
rect -61 -2208 -57 -2182
rect -10 -2191 -6 -2175
rect 17 -2177 21 -2167
rect 29 -2110 38 -2106
rect 91 -2107 95 -2103
rect 118 -2106 122 -2100
rect -20 -2194 -6 -2191
rect 29 -2192 32 -2110
rect 113 -2110 122 -2106
rect 42 -2118 56 -2114
rect 53 -2167 56 -2118
rect 42 -2171 56 -2167
rect 42 -2179 48 -2175
rect -61 -2212 -52 -2208
rect -61 -2233 -57 -2212
rect -48 -2220 -42 -2216
rect -61 -2237 -52 -2233
rect -61 -2252 -57 -2237
rect -45 -2241 -42 -2220
rect -27 -2234 -23 -2202
rect -20 -2209 -16 -2194
rect 29 -2196 38 -2192
rect 5 -2208 9 -2207
rect 0 -2212 9 -2208
rect -8 -2233 0 -2220
rect -48 -2245 -8 -2241
rect -61 -2255 -48 -2252
rect -48 -2258 -44 -2255
rect -48 -2262 -39 -2258
rect -22 -2259 -18 -2245
rect 5 -2258 9 -2212
rect 38 -2217 42 -2204
rect 38 -2225 42 -2222
rect 28 -2229 42 -2225
rect 28 -2252 31 -2229
rect 38 -2242 42 -2229
rect 45 -2250 48 -2179
rect 17 -2255 31 -2252
rect 42 -2254 48 -2250
rect 0 -2262 9 -2258
rect -35 -2270 -8 -2266
rect -22 -2278 -18 -2270
rect 5 -2277 9 -2262
rect 53 -2264 56 -2171
rect 59 -2118 105 -2114
rect 59 -2250 62 -2118
rect 118 -2125 122 -2115
rect 126 -2129 129 -2097
rect 91 -2132 129 -2129
rect 65 -2142 69 -2136
rect 65 -2146 74 -2142
rect 91 -2143 95 -2132
rect 118 -2142 122 -2141
rect 65 -2216 69 -2146
rect 113 -2146 122 -2142
rect 78 -2154 105 -2150
rect 91 -2168 95 -2154
rect 118 -2167 122 -2146
rect 113 -2171 122 -2167
rect 88 -2189 95 -2186
rect 85 -2211 88 -2191
rect 91 -2193 95 -2189
rect 105 -2192 113 -2179
rect 118 -2186 122 -2171
rect 113 -2204 128 -2200
rect 85 -2214 95 -2211
rect 70 -2217 78 -2216
rect 70 -2221 74 -2217
rect 91 -2218 95 -2214
rect 117 -2217 122 -2216
rect 65 -2236 69 -2221
rect 113 -2221 122 -2217
rect 78 -2229 105 -2225
rect 91 -2243 95 -2229
rect 118 -2236 122 -2221
rect 125 -2242 128 -2204
rect 113 -2246 128 -2242
rect 59 -2254 105 -2250
rect 125 -2264 128 -2246
rect 53 -2267 128 -2264
rect -73 -2281 -18 -2278
rect 125 -2359 128 -2267
rect 138 -2295 141 -2073
rect 148 -2274 152 -1906
rect 159 -1922 163 -1880
rect 284 -1883 287 -1862
rect 176 -1900 299 -1897
rect 159 -1926 168 -1922
rect 159 -1972 163 -1926
rect 168 -1947 172 -1934
rect 176 -1948 180 -1900
rect 295 -1903 299 -1900
rect 330 -1903 333 -1821
rect 439 -1832 443 -1791
rect 466 -1798 470 -1783
rect 514 -1785 517 -1692
rect 520 -1639 566 -1635
rect 520 -1771 523 -1639
rect 579 -1646 583 -1636
rect 587 -1650 590 -1618
rect 552 -1653 590 -1650
rect 526 -1663 530 -1657
rect 526 -1667 535 -1663
rect 552 -1664 556 -1653
rect 579 -1663 583 -1662
rect 526 -1737 530 -1667
rect 574 -1667 583 -1663
rect 539 -1675 566 -1671
rect 552 -1689 556 -1675
rect 579 -1688 583 -1667
rect 574 -1692 583 -1688
rect 549 -1710 556 -1707
rect 546 -1732 549 -1712
rect 552 -1714 556 -1710
rect 566 -1713 574 -1700
rect 579 -1707 583 -1692
rect 574 -1725 589 -1721
rect 546 -1735 556 -1732
rect 531 -1738 539 -1737
rect 531 -1742 535 -1738
rect 552 -1739 556 -1735
rect 578 -1738 583 -1737
rect 526 -1757 530 -1742
rect 574 -1742 583 -1738
rect 539 -1750 566 -1746
rect 552 -1764 556 -1750
rect 579 -1757 583 -1742
rect 586 -1763 589 -1725
rect 574 -1767 589 -1763
rect 520 -1775 566 -1771
rect 586 -1785 589 -1767
rect 514 -1788 589 -1785
rect 586 -1815 589 -1788
rect 605 -1822 608 -1365
rect 621 -1440 625 -1401
rect 740 -1406 743 -1032
rect 752 -1038 816 -1035
rect 638 -1418 755 -1415
rect 621 -1444 630 -1440
rect 621 -1490 625 -1444
rect 630 -1465 634 -1452
rect 638 -1466 642 -1418
rect 757 -1421 761 -1418
rect 923 -1419 926 -1032
rect 647 -1441 651 -1426
rect 757 -1424 795 -1421
rect 674 -1440 678 -1434
rect 669 -1444 678 -1440
rect 661 -1456 669 -1452
rect 647 -1461 669 -1456
rect 647 -1473 651 -1461
rect 661 -1465 669 -1461
rect 674 -1473 678 -1444
rect 634 -1477 651 -1473
rect 669 -1477 678 -1473
rect 621 -1494 630 -1490
rect 647 -1491 651 -1477
rect 674 -1490 678 -1477
rect 621 -1555 625 -1494
rect 669 -1494 678 -1490
rect 634 -1502 646 -1498
rect 651 -1502 661 -1498
rect 674 -1504 678 -1494
rect 695 -1437 704 -1433
rect 757 -1434 761 -1424
rect 784 -1433 788 -1427
rect 695 -1519 698 -1437
rect 779 -1437 788 -1433
rect 708 -1445 722 -1441
rect 719 -1494 722 -1445
rect 708 -1498 722 -1494
rect 708 -1506 714 -1502
rect 695 -1523 704 -1519
rect 704 -1544 708 -1531
rect 704 -1555 708 -1549
rect 621 -1560 708 -1555
rect 664 -1631 668 -1560
rect 704 -1569 708 -1560
rect 711 -1577 714 -1506
rect 708 -1581 714 -1577
rect 719 -1591 722 -1498
rect 725 -1445 771 -1441
rect 725 -1577 728 -1445
rect 784 -1452 788 -1442
rect 792 -1456 795 -1424
rect 757 -1459 795 -1456
rect 731 -1469 735 -1463
rect 731 -1473 740 -1469
rect 757 -1470 761 -1459
rect 784 -1469 788 -1468
rect 731 -1543 735 -1473
rect 779 -1473 788 -1469
rect 744 -1481 771 -1477
rect 757 -1495 761 -1481
rect 784 -1494 788 -1473
rect 779 -1498 788 -1494
rect 754 -1516 761 -1513
rect 751 -1538 754 -1518
rect 757 -1520 761 -1516
rect 771 -1519 779 -1506
rect 784 -1513 788 -1498
rect 779 -1531 794 -1527
rect 751 -1541 761 -1538
rect 736 -1548 740 -1544
rect 757 -1545 761 -1541
rect 783 -1544 788 -1543
rect 731 -1563 735 -1548
rect 779 -1548 788 -1544
rect 744 -1556 771 -1552
rect 757 -1570 761 -1556
rect 784 -1563 788 -1548
rect 791 -1569 794 -1531
rect 779 -1573 794 -1569
rect 725 -1581 771 -1577
rect 791 -1591 794 -1573
rect 719 -1594 794 -1591
rect 791 -1612 794 -1594
rect 804 -1604 808 -1419
rect 791 -1615 829 -1612
rect 791 -1618 795 -1615
rect 690 -1621 795 -1618
rect 664 -1635 673 -1631
rect 664 -1681 668 -1635
rect 673 -1656 677 -1643
rect 681 -1657 685 -1624
rect 690 -1632 694 -1621
rect 717 -1631 721 -1625
rect 712 -1635 721 -1631
rect 704 -1647 712 -1643
rect 690 -1652 712 -1647
rect 690 -1664 694 -1652
rect 704 -1656 712 -1652
rect 717 -1664 721 -1635
rect 677 -1668 694 -1664
rect 712 -1668 721 -1664
rect 664 -1685 673 -1681
rect 690 -1682 694 -1668
rect 717 -1681 721 -1668
rect 664 -1697 668 -1685
rect 712 -1685 721 -1681
rect 677 -1693 704 -1689
rect 639 -1700 668 -1697
rect 639 -1726 643 -1700
rect 690 -1709 694 -1693
rect 717 -1695 721 -1685
rect 729 -1628 738 -1624
rect 791 -1625 795 -1621
rect 818 -1624 822 -1618
rect 680 -1712 694 -1709
rect 729 -1710 732 -1628
rect 813 -1628 822 -1624
rect 742 -1636 756 -1632
rect 753 -1685 756 -1636
rect 742 -1689 756 -1685
rect 742 -1697 748 -1693
rect 639 -1730 648 -1726
rect 639 -1751 643 -1730
rect 652 -1738 658 -1734
rect 639 -1755 648 -1751
rect 639 -1770 643 -1755
rect 655 -1759 658 -1738
rect 673 -1752 677 -1720
rect 680 -1727 684 -1712
rect 729 -1714 738 -1710
rect 705 -1726 709 -1725
rect 700 -1730 709 -1726
rect 692 -1751 700 -1738
rect 652 -1763 692 -1759
rect 639 -1773 652 -1770
rect 652 -1776 656 -1773
rect 652 -1780 661 -1776
rect 678 -1777 682 -1763
rect 705 -1776 709 -1730
rect 738 -1735 742 -1722
rect 738 -1743 742 -1740
rect 728 -1747 742 -1743
rect 728 -1770 731 -1747
rect 738 -1760 742 -1747
rect 745 -1768 748 -1697
rect 717 -1773 731 -1770
rect 742 -1772 748 -1768
rect 652 -1795 656 -1780
rect 700 -1780 709 -1776
rect 665 -1788 692 -1784
rect 678 -1805 682 -1788
rect 705 -1795 709 -1780
rect 753 -1782 756 -1689
rect 759 -1636 805 -1632
rect 759 -1768 762 -1636
rect 818 -1643 822 -1633
rect 826 -1647 829 -1615
rect 791 -1650 829 -1647
rect 765 -1660 769 -1654
rect 765 -1664 774 -1660
rect 791 -1661 795 -1650
rect 818 -1660 822 -1659
rect 765 -1734 769 -1664
rect 813 -1664 822 -1660
rect 778 -1672 805 -1668
rect 791 -1686 795 -1672
rect 818 -1685 822 -1664
rect 813 -1689 822 -1685
rect 788 -1707 795 -1704
rect 785 -1729 788 -1709
rect 791 -1711 795 -1707
rect 805 -1710 813 -1697
rect 818 -1704 822 -1689
rect 813 -1722 828 -1718
rect 785 -1732 795 -1729
rect 770 -1735 778 -1734
rect 770 -1739 774 -1735
rect 791 -1736 795 -1732
rect 817 -1735 822 -1734
rect 765 -1754 769 -1739
rect 813 -1739 822 -1735
rect 778 -1747 805 -1743
rect 791 -1761 795 -1747
rect 818 -1754 822 -1739
rect 825 -1760 828 -1722
rect 813 -1764 828 -1760
rect 759 -1772 805 -1768
rect 825 -1782 828 -1764
rect 753 -1785 828 -1782
rect 605 -1825 718 -1822
rect 295 -1906 333 -1903
rect 185 -1923 189 -1908
rect 212 -1922 216 -1916
rect 207 -1926 216 -1922
rect 199 -1938 207 -1934
rect 185 -1943 207 -1938
rect 185 -1955 189 -1943
rect 199 -1947 207 -1943
rect 212 -1955 216 -1926
rect 172 -1959 189 -1955
rect 207 -1959 216 -1955
rect 159 -1976 168 -1972
rect 185 -1973 189 -1959
rect 212 -1972 216 -1959
rect 159 -2037 163 -1976
rect 207 -1976 216 -1972
rect 172 -1984 184 -1980
rect 189 -1984 199 -1980
rect 212 -1986 216 -1976
rect 233 -1919 242 -1915
rect 295 -1916 299 -1906
rect 322 -1915 326 -1909
rect 233 -2001 236 -1919
rect 317 -1919 326 -1915
rect 246 -1927 260 -1923
rect 257 -1976 260 -1927
rect 246 -1980 260 -1976
rect 246 -1988 252 -1984
rect 233 -2005 242 -2001
rect 242 -2026 246 -2013
rect 242 -2037 246 -2031
rect 159 -2042 246 -2037
rect 202 -2113 206 -2042
rect 242 -2051 246 -2042
rect 249 -2059 252 -1988
rect 246 -2063 252 -2059
rect 257 -2073 260 -1980
rect 263 -1927 309 -1923
rect 263 -2059 266 -1927
rect 322 -1934 326 -1924
rect 330 -1938 333 -1906
rect 295 -1941 333 -1938
rect 342 -1835 443 -1832
rect 269 -1951 273 -1945
rect 269 -1955 278 -1951
rect 295 -1952 299 -1941
rect 322 -1951 326 -1950
rect 269 -2025 273 -1955
rect 317 -1955 326 -1951
rect 282 -1963 309 -1959
rect 295 -1977 299 -1963
rect 322 -1976 326 -1955
rect 317 -1980 326 -1976
rect 292 -1998 299 -1995
rect 289 -2020 292 -2000
rect 295 -2002 299 -1998
rect 309 -2001 317 -1988
rect 322 -1995 326 -1980
rect 317 -2013 332 -2009
rect 289 -2023 299 -2020
rect 274 -2030 278 -2026
rect 295 -2027 299 -2023
rect 321 -2026 326 -2025
rect 269 -2045 273 -2030
rect 317 -2030 326 -2026
rect 282 -2038 309 -2034
rect 295 -2052 299 -2038
rect 322 -2045 326 -2030
rect 329 -2051 332 -2013
rect 317 -2055 332 -2051
rect 263 -2063 309 -2059
rect 329 -2073 332 -2055
rect 257 -2076 332 -2073
rect 329 -2094 332 -2076
rect 342 -2086 346 -1835
rect 376 -1871 526 -1868
rect 329 -2097 367 -2094
rect 329 -2100 333 -2097
rect 228 -2103 333 -2100
rect 202 -2117 211 -2113
rect 202 -2163 206 -2117
rect 211 -2138 215 -2125
rect 219 -2139 223 -2106
rect 228 -2114 232 -2103
rect 255 -2113 259 -2107
rect 250 -2117 259 -2113
rect 242 -2129 250 -2125
rect 228 -2134 250 -2129
rect 228 -2146 232 -2134
rect 242 -2138 250 -2134
rect 255 -2146 259 -2117
rect 215 -2150 232 -2146
rect 250 -2150 259 -2146
rect 202 -2167 211 -2163
rect 228 -2164 232 -2150
rect 255 -2163 259 -2150
rect 202 -2179 206 -2167
rect 250 -2167 259 -2163
rect 215 -2175 242 -2171
rect 177 -2182 206 -2179
rect 177 -2208 181 -2182
rect 228 -2191 232 -2175
rect 255 -2177 259 -2167
rect 267 -2110 276 -2106
rect 329 -2107 333 -2103
rect 356 -2106 360 -2100
rect 218 -2194 232 -2191
rect 267 -2192 270 -2110
rect 351 -2110 360 -2106
rect 280 -2118 294 -2114
rect 291 -2167 294 -2118
rect 280 -2171 294 -2167
rect 280 -2179 286 -2175
rect 177 -2212 186 -2208
rect 177 -2233 181 -2212
rect 190 -2220 196 -2216
rect 177 -2237 186 -2233
rect 177 -2252 181 -2237
rect 193 -2241 196 -2220
rect 211 -2234 215 -2202
rect 218 -2209 222 -2194
rect 267 -2196 276 -2192
rect 243 -2208 247 -2207
rect 238 -2212 247 -2208
rect 230 -2233 238 -2220
rect 190 -2245 230 -2241
rect 177 -2255 190 -2252
rect 190 -2258 194 -2255
rect 190 -2262 199 -2258
rect 216 -2259 220 -2245
rect 243 -2258 247 -2212
rect 276 -2217 280 -2204
rect 276 -2225 280 -2222
rect 266 -2229 280 -2225
rect 266 -2252 269 -2229
rect 276 -2242 280 -2229
rect 283 -2250 286 -2179
rect 255 -2255 269 -2252
rect 280 -2254 286 -2250
rect 238 -2262 247 -2258
rect 203 -2270 230 -2266
rect 216 -2274 220 -2270
rect 148 -2277 220 -2274
rect 243 -2277 247 -2262
rect 291 -2264 294 -2171
rect 297 -2118 343 -2114
rect 297 -2250 300 -2118
rect 356 -2125 360 -2115
rect 364 -2129 367 -2097
rect 329 -2132 367 -2129
rect 303 -2142 307 -2136
rect 303 -2146 312 -2142
rect 329 -2143 333 -2132
rect 356 -2142 360 -2141
rect 303 -2216 307 -2146
rect 351 -2146 360 -2142
rect 316 -2154 343 -2150
rect 329 -2168 333 -2154
rect 356 -2167 360 -2146
rect 351 -2171 360 -2167
rect 326 -2189 333 -2186
rect 323 -2211 326 -2191
rect 329 -2193 333 -2189
rect 343 -2192 351 -2179
rect 356 -2186 360 -2171
rect 351 -2204 366 -2200
rect 323 -2214 333 -2211
rect 308 -2217 316 -2216
rect 308 -2221 312 -2217
rect 329 -2218 333 -2214
rect 355 -2217 360 -2216
rect 303 -2236 307 -2221
rect 351 -2221 360 -2217
rect 316 -2229 343 -2225
rect 329 -2243 333 -2229
rect 356 -2236 360 -2221
rect 363 -2242 366 -2204
rect 351 -2246 366 -2242
rect 297 -2254 343 -2250
rect 363 -2264 366 -2246
rect 291 -2267 366 -2264
rect 363 -2288 366 -2267
rect 376 -2288 379 -1871
rect 403 -1911 407 -1880
rect 420 -1889 543 -1886
rect 403 -1915 412 -1911
rect 403 -1961 407 -1915
rect 412 -1936 416 -1923
rect 420 -1937 424 -1889
rect 539 -1892 543 -1889
rect 539 -1895 590 -1892
rect 429 -1912 433 -1897
rect 456 -1911 460 -1905
rect 451 -1915 460 -1911
rect 443 -1927 451 -1923
rect 429 -1932 451 -1927
rect 429 -1944 433 -1932
rect 443 -1936 451 -1932
rect 456 -1944 460 -1915
rect 416 -1948 433 -1944
rect 451 -1948 460 -1944
rect 403 -1965 412 -1961
rect 429 -1962 433 -1948
rect 456 -1961 460 -1948
rect 403 -2007 407 -1965
rect 451 -1965 460 -1961
rect 416 -1973 428 -1969
rect 433 -1973 443 -1969
rect 456 -1975 460 -1965
rect 477 -1908 486 -1904
rect 539 -1905 543 -1895
rect 566 -1904 570 -1898
rect 477 -1990 480 -1908
rect 561 -1908 570 -1904
rect 490 -1916 504 -1912
rect 501 -1965 504 -1916
rect 490 -1969 504 -1965
rect 490 -1977 496 -1973
rect 477 -1994 486 -1990
rect 486 -2007 490 -2002
rect 403 -2012 490 -2007
rect 486 -2015 490 -2012
rect 486 -2040 490 -2020
rect 493 -2048 496 -1977
rect 490 -2052 496 -2048
rect 501 -2062 504 -1969
rect 507 -1916 553 -1912
rect 507 -2048 510 -1916
rect 566 -1923 570 -1913
rect 574 -1927 577 -1895
rect 539 -1930 577 -1927
rect 513 -1940 517 -1934
rect 513 -1944 522 -1940
rect 539 -1941 543 -1930
rect 566 -1940 570 -1939
rect 513 -2014 517 -1944
rect 561 -1944 570 -1940
rect 526 -1952 553 -1948
rect 539 -1966 543 -1952
rect 566 -1965 570 -1944
rect 561 -1969 570 -1965
rect 536 -1987 543 -1984
rect 533 -2009 536 -1989
rect 539 -1991 543 -1987
rect 553 -1990 561 -1977
rect 566 -1984 570 -1969
rect 561 -2002 576 -1998
rect 533 -2012 543 -2009
rect 518 -2019 522 -2015
rect 539 -2016 543 -2012
rect 565 -2015 570 -2014
rect 513 -2034 517 -2019
rect 561 -2019 570 -2015
rect 526 -2027 553 -2023
rect 539 -2041 543 -2027
rect 566 -2034 570 -2019
rect 573 -2040 576 -2002
rect 561 -2044 576 -2040
rect 507 -2052 553 -2048
rect 573 -2062 576 -2044
rect 501 -2065 576 -2062
rect 363 -2291 379 -2288
rect 429 -2295 433 -2135
rect 138 -2298 433 -2295
rect 573 -2359 576 -2065
rect 587 -2270 590 -1895
rect 596 -1919 600 -1880
rect 715 -1885 718 -1825
rect 613 -1897 730 -1894
rect 596 -1923 605 -1919
rect 596 -1969 600 -1923
rect 605 -1944 609 -1931
rect 613 -1945 617 -1897
rect 732 -1900 736 -1897
rect 732 -1903 770 -1900
rect 622 -1920 626 -1905
rect 649 -1919 653 -1913
rect 644 -1923 653 -1919
rect 636 -1935 644 -1931
rect 622 -1940 644 -1935
rect 622 -1952 626 -1940
rect 636 -1944 644 -1940
rect 649 -1952 653 -1923
rect 609 -1956 626 -1952
rect 644 -1956 653 -1952
rect 596 -1973 605 -1969
rect 622 -1970 626 -1956
rect 649 -1969 653 -1956
rect 596 -2034 600 -1973
rect 644 -1973 653 -1969
rect 609 -1981 621 -1977
rect 626 -1981 636 -1977
rect 649 -1983 653 -1973
rect 670 -1916 679 -1912
rect 732 -1913 736 -1903
rect 759 -1912 763 -1906
rect 670 -1998 673 -1916
rect 754 -1916 763 -1912
rect 683 -1924 697 -1920
rect 694 -1973 697 -1924
rect 683 -1977 697 -1973
rect 683 -1985 689 -1981
rect 670 -2002 679 -1998
rect 679 -2023 683 -2010
rect 679 -2034 683 -2028
rect 596 -2039 683 -2034
rect 639 -2110 643 -2039
rect 679 -2048 683 -2039
rect 686 -2056 689 -1985
rect 683 -2060 689 -2056
rect 694 -2070 697 -1977
rect 700 -1924 746 -1920
rect 700 -2056 703 -1924
rect 759 -1931 763 -1921
rect 767 -1935 770 -1903
rect 732 -1938 770 -1935
rect 706 -1948 710 -1942
rect 706 -1952 715 -1948
rect 732 -1949 736 -1938
rect 759 -1948 763 -1947
rect 706 -2022 710 -1952
rect 754 -1952 763 -1948
rect 719 -1960 746 -1956
rect 732 -1974 736 -1960
rect 759 -1973 763 -1952
rect 754 -1977 763 -1973
rect 729 -1995 736 -1992
rect 726 -2017 729 -1997
rect 732 -1999 736 -1995
rect 746 -1998 754 -1985
rect 759 -1992 763 -1977
rect 754 -2010 769 -2006
rect 726 -2020 736 -2017
rect 711 -2027 715 -2023
rect 732 -2024 736 -2020
rect 758 -2023 763 -2022
rect 706 -2042 710 -2027
rect 754 -2027 763 -2023
rect 719 -2035 746 -2031
rect 732 -2049 736 -2035
rect 759 -2042 763 -2027
rect 766 -2048 769 -2010
rect 754 -2052 769 -2048
rect 700 -2060 746 -2056
rect 766 -2070 769 -2052
rect 694 -2073 769 -2070
rect 766 -2091 769 -2073
rect 779 -2083 783 -1898
rect 766 -2094 804 -2091
rect 766 -2097 770 -2094
rect 665 -2100 770 -2097
rect 639 -2114 648 -2110
rect 639 -2160 643 -2114
rect 648 -2135 652 -2122
rect 656 -2136 660 -2103
rect 665 -2111 669 -2100
rect 692 -2110 696 -2104
rect 687 -2114 696 -2110
rect 679 -2126 687 -2122
rect 665 -2131 687 -2126
rect 665 -2143 669 -2131
rect 679 -2135 687 -2131
rect 692 -2143 696 -2114
rect 652 -2147 669 -2143
rect 687 -2147 696 -2143
rect 639 -2164 648 -2160
rect 665 -2161 669 -2147
rect 692 -2160 696 -2147
rect 639 -2176 643 -2164
rect 687 -2164 696 -2160
rect 652 -2172 679 -2168
rect 614 -2179 643 -2176
rect 614 -2205 618 -2179
rect 665 -2188 669 -2172
rect 692 -2174 696 -2164
rect 704 -2107 713 -2103
rect 766 -2104 770 -2100
rect 793 -2103 797 -2097
rect 655 -2191 669 -2188
rect 704 -2189 707 -2107
rect 788 -2107 797 -2103
rect 717 -2115 731 -2111
rect 728 -2164 731 -2115
rect 717 -2168 731 -2164
rect 717 -2176 723 -2172
rect 614 -2209 623 -2205
rect 614 -2230 618 -2209
rect 627 -2217 633 -2213
rect 614 -2234 623 -2230
rect 614 -2249 618 -2234
rect 630 -2238 633 -2217
rect 648 -2231 652 -2199
rect 655 -2206 659 -2191
rect 704 -2193 713 -2189
rect 680 -2205 684 -2204
rect 675 -2209 684 -2205
rect 667 -2230 675 -2217
rect 627 -2242 667 -2238
rect 614 -2252 627 -2249
rect 627 -2255 631 -2252
rect 627 -2259 636 -2255
rect 653 -2256 657 -2242
rect 680 -2255 684 -2209
rect 713 -2214 717 -2201
rect 713 -2222 717 -2219
rect 703 -2226 717 -2222
rect 703 -2249 706 -2226
rect 713 -2239 717 -2226
rect 720 -2247 723 -2176
rect 692 -2252 706 -2249
rect 717 -2251 723 -2247
rect 675 -2259 684 -2255
rect 640 -2267 667 -2263
rect 653 -2270 657 -2267
rect 587 -2274 657 -2270
rect 680 -2274 684 -2259
rect 728 -2261 731 -2168
rect 734 -2115 780 -2111
rect 734 -2247 737 -2115
rect 793 -2122 797 -2112
rect 801 -2126 804 -2094
rect 766 -2129 804 -2126
rect 740 -2139 744 -2133
rect 740 -2143 749 -2139
rect 766 -2140 770 -2129
rect 793 -2139 797 -2138
rect 740 -2213 744 -2143
rect 788 -2143 797 -2139
rect 753 -2151 780 -2147
rect 766 -2165 770 -2151
rect 793 -2164 797 -2143
rect 788 -2168 797 -2164
rect 763 -2186 770 -2183
rect 760 -2208 763 -2188
rect 766 -2190 770 -2186
rect 780 -2189 788 -2176
rect 793 -2183 797 -2168
rect 788 -2201 803 -2197
rect 760 -2211 770 -2208
rect 745 -2214 753 -2213
rect 745 -2218 749 -2214
rect 766 -2215 770 -2211
rect 792 -2214 797 -2213
rect 740 -2233 744 -2218
rect 788 -2218 797 -2214
rect 753 -2226 780 -2222
rect 766 -2240 770 -2226
rect 793 -2233 797 -2218
rect 800 -2239 803 -2201
rect 788 -2243 803 -2239
rect 734 -2251 780 -2247
rect 800 -2261 803 -2243
rect 728 -2264 803 -2261
rect 800 -2358 803 -2264
rect 825 -2357 828 -1785
rect 923 -2356 927 -1419
rect 937 -2356 941 -816
rect 964 -823 968 -808
rect 994 -1032 999 -745
rect 994 -1796 999 -1038
rect 994 -2275 999 -1801
<< m2contact >>
rect 36 -680 41 -675
rect 96 -680 101 -675
rect 276 -680 281 -675
rect 456 -680 461 -675
rect 156 -688 161 -683
rect 336 -688 341 -683
rect 396 -688 401 -683
rect 696 -688 701 -683
rect 216 -696 221 -691
rect 576 -696 581 -691
rect 636 -696 641 -691
rect 816 -696 821 -691
rect 516 -704 521 -699
rect 756 -704 761 -699
rect 876 -704 881 -699
rect 927 -704 932 -699
rect 28 -714 33 -709
rect 147 -714 152 -709
rect 207 -714 212 -709
rect 507 -714 512 -709
rect 87 -722 92 -717
rect 327 -722 332 -717
rect 567 -722 572 -717
rect 747 -722 752 -717
rect 267 -730 272 -725
rect 387 -730 392 -725
rect 627 -730 632 -725
rect 867 -730 872 -725
rect 447 -738 452 -733
rect 687 -738 692 -733
rect 807 -738 812 -733
rect 936 -738 941 -733
rect 27 -753 32 -748
rect 36 -752 41 -747
rect 10 -830 15 -825
rect 87 -753 92 -748
rect 96 -752 101 -747
rect 70 -831 75 -826
rect -276 -1402 -270 -1397
rect 147 -753 152 -748
rect 156 -752 161 -747
rect 130 -831 135 -826
rect 207 -753 212 -748
rect 216 -752 221 -747
rect 190 -831 195 -826
rect 112 -864 118 -859
rect 14 -880 19 -875
rect 13 -957 18 -952
rect 41 -963 46 -958
rect 70 -1003 75 -998
rect 151 -896 156 -891
rect 151 -922 156 -917
rect 116 -972 121 -967
rect 98 -1002 103 -997
rect 150 -997 155 -992
rect 171 -1063 176 -1058
rect 48 -1078 53 -1073
rect 84 -1154 89 -1149
rect 39 -1174 44 -1169
rect 72 -1179 77 -1174
rect 19 -1227 24 -1222
rect 104 -1194 109 -1189
rect 79 -1227 84 -1222
rect 17 -1262 23 -1256
rect 185 -1087 190 -1082
rect 185 -1113 190 -1108
rect 150 -1163 155 -1158
rect 132 -1193 137 -1188
rect 184 -1188 189 -1183
rect 126 -1280 132 -1274
rect -250 -1430 -245 -1425
rect -251 -1507 -246 -1502
rect -223 -1513 -218 -1508
rect -194 -1553 -189 -1548
rect -113 -1446 -108 -1441
rect -113 -1472 -108 -1467
rect -148 -1522 -143 -1517
rect -166 -1552 -161 -1547
rect -114 -1547 -109 -1542
rect -93 -1613 -88 -1608
rect -216 -1628 -211 -1623
rect -180 -1704 -175 -1699
rect -225 -1724 -220 -1719
rect -192 -1729 -187 -1724
rect -245 -1777 -240 -1772
rect -160 -1744 -155 -1739
rect -185 -1777 -180 -1772
rect -79 -1637 -74 -1632
rect -79 -1663 -74 -1658
rect -114 -1713 -109 -1708
rect -132 -1743 -127 -1738
rect -80 -1738 -75 -1733
rect -79 -1880 -73 -1875
rect 267 -753 272 -748
rect 276 -752 281 -747
rect 250 -831 255 -826
rect 327 -753 332 -748
rect 336 -752 341 -747
rect 310 -831 315 -826
rect 387 -753 392 -748
rect 396 -752 401 -747
rect 370 -831 375 -826
rect 447 -753 452 -748
rect 456 -752 461 -747
rect 430 -831 435 -826
rect 396 -840 401 -835
rect 507 -753 512 -748
rect 516 -752 521 -747
rect 490 -831 495 -826
rect 567 -753 572 -748
rect 576 -752 581 -747
rect 550 -831 555 -826
rect 627 -753 632 -748
rect 636 -752 641 -747
rect 610 -831 615 -826
rect 687 -753 692 -748
rect 696 -752 701 -747
rect 670 -831 675 -826
rect 747 -753 752 -748
rect 756 -752 761 -747
rect 730 -831 735 -826
rect 807 -753 812 -748
rect 816 -752 821 -747
rect 790 -831 795 -826
rect 633 -844 638 -839
rect 867 -753 872 -748
rect 876 -752 881 -747
rect 850 -831 855 -826
rect 816 -845 821 -840
rect 927 -753 932 -748
rect 936 -752 941 -747
rect 910 -831 915 -826
rect 217 -1282 222 -1276
rect 153 -1401 159 -1396
rect 359 -860 364 -855
rect 358 -937 363 -932
rect 386 -943 391 -938
rect 373 -975 379 -970
rect 415 -983 420 -978
rect 334 -991 340 -986
rect 179 -1429 184 -1424
rect 178 -1506 183 -1501
rect 206 -1512 211 -1507
rect 235 -1552 240 -1547
rect 316 -1445 321 -1440
rect 316 -1471 321 -1466
rect 281 -1521 286 -1516
rect 263 -1551 268 -1546
rect 315 -1546 320 -1541
rect 496 -876 501 -871
rect 496 -902 501 -897
rect 461 -952 466 -947
rect 596 -864 601 -859
rect 443 -982 448 -977
rect 495 -977 500 -972
rect 595 -941 600 -936
rect 623 -947 628 -942
rect 607 -979 612 -974
rect 652 -987 657 -982
rect 360 -1036 366 -1029
rect 396 -1036 402 -1029
rect 382 -1401 388 -1396
rect 733 -880 738 -875
rect 733 -906 738 -901
rect 698 -956 703 -951
rect 779 -864 784 -859
rect 680 -986 685 -981
rect 732 -981 737 -976
rect 778 -941 783 -936
rect 806 -947 811 -942
rect 794 -979 799 -974
rect 835 -987 840 -982
rect 510 -1038 516 -1031
rect 632 -1038 638 -1031
rect 916 -880 921 -875
rect 916 -906 921 -901
rect 881 -956 886 -951
rect 863 -986 868 -981
rect 915 -981 920 -976
rect 408 -1429 413 -1424
rect 407 -1506 412 -1501
rect 435 -1512 440 -1507
rect 464 -1552 469 -1547
rect 336 -1612 341 -1607
rect 213 -1627 218 -1622
rect 249 -1703 254 -1698
rect 204 -1723 209 -1718
rect 237 -1728 242 -1723
rect 184 -1776 189 -1771
rect 269 -1743 274 -1738
rect 244 -1776 249 -1771
rect 350 -1636 355 -1631
rect 545 -1445 550 -1440
rect 545 -1471 550 -1466
rect 510 -1521 515 -1516
rect 492 -1551 497 -1546
rect 544 -1546 549 -1541
rect 565 -1612 570 -1607
rect 442 -1627 447 -1622
rect 350 -1662 355 -1657
rect 315 -1712 320 -1707
rect 297 -1742 302 -1737
rect 349 -1737 354 -1732
rect 478 -1703 483 -1698
rect 433 -1723 438 -1718
rect 466 -1728 471 -1723
rect 413 -1776 418 -1771
rect 498 -1743 503 -1738
rect 473 -1776 478 -1771
rect 159 -1880 165 -1875
rect 44 -1888 51 -1883
rect -53 -1908 -48 -1903
rect -54 -1985 -49 -1980
rect -26 -1991 -21 -1986
rect 3 -2031 8 -2026
rect 84 -1924 89 -1919
rect 84 -1950 89 -1945
rect 49 -2000 54 -1995
rect 31 -2030 36 -2025
rect 83 -2025 88 -2020
rect 104 -2091 109 -2086
rect -19 -2106 -14 -2101
rect 17 -2182 22 -2177
rect -28 -2202 -23 -2197
rect 5 -2207 10 -2202
rect -48 -2255 -43 -2250
rect 37 -2222 42 -2217
rect 12 -2255 17 -2250
rect 118 -2115 123 -2110
rect 118 -2141 123 -2136
rect 83 -2191 88 -2186
rect 65 -2221 70 -2216
rect 117 -2216 122 -2211
rect 282 -1888 289 -1883
rect 579 -1636 584 -1631
rect 579 -1662 584 -1657
rect 544 -1712 549 -1707
rect 526 -1742 531 -1737
rect 578 -1737 583 -1732
rect 621 -1401 627 -1396
rect 747 -1040 752 -1035
rect 816 -1040 821 -1035
rect 647 -1426 652 -1421
rect 646 -1503 651 -1498
rect 674 -1509 679 -1504
rect 703 -1549 708 -1544
rect 784 -1442 789 -1437
rect 784 -1468 789 -1463
rect 749 -1518 754 -1513
rect 731 -1548 736 -1543
rect 783 -1543 788 -1538
rect 804 -1609 809 -1604
rect 681 -1624 686 -1619
rect 717 -1700 722 -1695
rect 672 -1720 677 -1715
rect 705 -1725 710 -1720
rect 652 -1773 657 -1768
rect 737 -1740 742 -1735
rect 712 -1773 717 -1768
rect 818 -1633 823 -1628
rect 818 -1659 823 -1654
rect 783 -1709 788 -1704
rect 765 -1739 770 -1734
rect 817 -1734 822 -1729
rect 185 -1908 190 -1903
rect 184 -1985 189 -1980
rect 212 -1991 217 -1986
rect 241 -2031 246 -2026
rect 322 -1924 327 -1919
rect 322 -1950 327 -1945
rect 287 -2000 292 -1995
rect 269 -2030 274 -2025
rect 321 -2025 326 -2020
rect 342 -2091 347 -2086
rect 219 -2106 224 -2101
rect 255 -2182 260 -2177
rect 210 -2202 215 -2197
rect 243 -2207 248 -2202
rect 190 -2255 195 -2250
rect 275 -2222 280 -2217
rect 250 -2255 255 -2250
rect 356 -2115 361 -2110
rect 356 -2141 361 -2136
rect 321 -2191 326 -2186
rect 303 -2221 308 -2216
rect 355 -2216 360 -2211
rect 403 -1880 409 -1875
rect 596 -1880 602 -1875
rect 429 -1897 434 -1892
rect 428 -1974 433 -1969
rect 456 -1980 461 -1975
rect 485 -2020 490 -2015
rect 566 -1913 571 -1908
rect 566 -1939 571 -1934
rect 531 -1989 536 -1984
rect 513 -2019 518 -2014
rect 565 -2014 570 -2009
rect 428 -2135 434 -2130
rect 622 -1905 627 -1900
rect 621 -1982 626 -1977
rect 649 -1988 654 -1983
rect 678 -2028 683 -2023
rect 759 -1921 764 -1916
rect 759 -1947 764 -1942
rect 724 -1997 729 -1992
rect 706 -2027 711 -2022
rect 758 -2022 763 -2017
rect 779 -2088 784 -2083
rect 656 -2103 661 -2098
rect 692 -2179 697 -2174
rect 647 -2199 652 -2194
rect 680 -2204 685 -2199
rect 627 -2252 632 -2247
rect 712 -2219 717 -2214
rect 687 -2252 692 -2247
rect 793 -2112 798 -2107
rect 793 -2138 798 -2133
rect 758 -2188 763 -2183
rect 740 -2218 745 -2213
rect 792 -2213 797 -2208
rect 994 -1038 999 -1032
rect 994 -1801 999 -1796
rect 992 -2282 1001 -2275
<< metal2 >>
rect 28 -748 32 -714
rect 37 -747 41 -680
rect 88 -748 92 -722
rect 97 -747 101 -680
rect 148 -748 152 -714
rect 157 -747 161 -688
rect 208 -748 212 -714
rect 217 -747 221 -696
rect 268 -748 272 -730
rect 277 -747 281 -680
rect 328 -748 332 -722
rect 337 -747 341 -688
rect 388 -748 392 -730
rect 397 -747 401 -688
rect 448 -748 452 -738
rect 457 -747 461 -680
rect 508 -748 512 -714
rect 517 -747 521 -704
rect 568 -748 572 -722
rect 577 -747 581 -696
rect 628 -748 632 -730
rect 637 -747 641 -696
rect 688 -748 692 -738
rect 697 -747 701 -688
rect 748 -748 752 -722
rect 757 -747 761 -704
rect 808 -748 812 -738
rect 817 -747 821 -696
rect 868 -748 872 -730
rect 877 -747 881 -704
rect 928 -748 932 -704
rect 937 -747 941 -738
rect -309 -830 10 -827
rect 15 -830 70 -827
rect -309 -1258 -305 -830
rect 75 -830 130 -827
rect 135 -830 190 -827
rect 195 -830 250 -827
rect 255 -830 310 -827
rect 315 -830 370 -827
rect 375 -830 430 -827
rect 435 -830 490 -827
rect 495 -830 550 -827
rect 555 -830 610 -827
rect 615 -830 670 -827
rect 675 -830 730 -827
rect 735 -830 790 -827
rect 795 -830 850 -827
rect 855 -830 910 -827
rect 397 -855 401 -840
rect 364 -858 461 -855
rect 113 -875 116 -864
rect 19 -878 116 -875
rect 14 -1162 18 -957
rect 46 -963 56 -958
rect 53 -1051 56 -963
rect 113 -972 116 -878
rect 156 -896 168 -891
rect 165 -917 168 -896
rect 156 -922 168 -917
rect 165 -992 168 -922
rect 359 -988 363 -937
rect 391 -943 401 -938
rect 340 -991 363 -988
rect 155 -997 168 -992
rect 75 -1002 98 -998
rect 165 -1031 168 -997
rect 165 -1034 360 -1031
rect 165 -1051 168 -1034
rect 375 -1046 379 -975
rect 398 -1029 401 -943
rect 458 -952 461 -858
rect 634 -859 638 -844
rect 817 -859 821 -845
rect 601 -862 698 -859
rect 501 -876 513 -871
rect 510 -897 513 -876
rect 501 -902 513 -897
rect 510 -972 513 -902
rect 500 -977 513 -972
rect 420 -982 443 -978
rect 510 -1031 513 -977
rect 596 -989 600 -941
rect 628 -947 638 -942
rect 402 -1034 510 -1031
rect 609 -1046 612 -979
rect 635 -1031 638 -947
rect 695 -956 698 -862
rect 784 -862 881 -859
rect 738 -880 750 -875
rect 747 -901 750 -880
rect 738 -906 750 -901
rect 747 -976 750 -906
rect 737 -981 750 -976
rect 657 -986 680 -982
rect 747 -1035 750 -981
rect 779 -993 783 -941
rect 811 -947 821 -942
rect 638 -1038 747 -1035
rect 796 -1046 799 -979
rect 818 -1035 821 -947
rect 878 -956 881 -862
rect 921 -880 933 -875
rect 930 -901 933 -880
rect 921 -906 933 -901
rect 930 -976 933 -906
rect 920 -981 933 -976
rect 840 -986 863 -982
rect 930 -1035 933 -981
rect 821 -1038 994 -1035
rect 237 -1049 799 -1046
rect 53 -1054 202 -1051
rect 147 -1063 171 -1060
rect 147 -1066 150 -1063
rect 48 -1069 150 -1066
rect 48 -1073 52 -1069
rect 14 -1165 44 -1162
rect 40 -1169 44 -1165
rect 89 -1174 92 -1149
rect 147 -1163 150 -1069
rect 199 -1082 202 -1054
rect 190 -1087 202 -1082
rect 199 -1108 202 -1087
rect 190 -1113 202 -1108
rect 77 -1178 92 -1174
rect 24 -1227 79 -1224
rect 89 -1242 92 -1178
rect 199 -1183 202 -1113
rect 189 -1188 202 -1183
rect 109 -1193 132 -1189
rect 199 -1242 202 -1188
rect 89 -1246 202 -1242
rect 199 -1248 202 -1246
rect -309 -1262 17 -1258
rect 23 -1262 139 -1258
rect -309 -1397 -305 -1262
rect 136 -1266 139 -1262
rect 237 -1266 241 -1049
rect 136 -1270 241 -1266
rect 132 -1279 217 -1276
rect 40 -1397 153 -1396
rect -309 -1400 -276 -1397
rect -309 -1875 -305 -1400
rect -270 -1399 153 -1397
rect -270 -1400 73 -1399
rect 159 -1399 382 -1396
rect 388 -1399 621 -1396
rect -245 -1428 -154 -1425
rect 184 -1427 275 -1424
rect 413 -1427 504 -1424
rect 652 -1424 743 -1421
rect -250 -1712 -246 -1507
rect -218 -1513 -208 -1508
rect -211 -1601 -208 -1513
rect -151 -1522 -148 -1431
rect -108 -1446 -96 -1441
rect -99 -1467 -96 -1446
rect -108 -1472 -96 -1467
rect -99 -1542 -96 -1472
rect -109 -1547 -96 -1542
rect -189 -1552 -166 -1548
rect -99 -1601 -96 -1547
rect -211 -1604 -62 -1601
rect -117 -1613 -93 -1610
rect -117 -1616 -114 -1613
rect -216 -1619 -114 -1616
rect -216 -1623 -212 -1619
rect -250 -1715 -220 -1712
rect -224 -1719 -220 -1715
rect -175 -1724 -172 -1699
rect -117 -1713 -114 -1619
rect -65 -1632 -62 -1604
rect -74 -1637 -62 -1632
rect -65 -1658 -62 -1637
rect -74 -1663 -62 -1658
rect -187 -1728 -172 -1724
rect -240 -1777 -185 -1774
rect -175 -1792 -172 -1728
rect -65 -1733 -62 -1663
rect 179 -1711 183 -1506
rect 211 -1512 221 -1507
rect 218 -1600 221 -1512
rect 278 -1521 281 -1430
rect 321 -1445 333 -1440
rect 330 -1466 333 -1445
rect 321 -1471 333 -1466
rect 330 -1541 333 -1471
rect 320 -1546 333 -1541
rect 240 -1551 263 -1547
rect 330 -1600 333 -1546
rect 218 -1603 367 -1600
rect 312 -1612 336 -1609
rect 312 -1615 315 -1612
rect 213 -1618 315 -1615
rect 213 -1622 217 -1618
rect 179 -1714 209 -1711
rect 205 -1718 209 -1714
rect 254 -1723 257 -1698
rect 312 -1712 315 -1618
rect 364 -1631 367 -1603
rect 355 -1636 367 -1631
rect 364 -1657 367 -1636
rect 355 -1662 367 -1657
rect 242 -1727 257 -1723
rect -75 -1738 -62 -1733
rect -155 -1743 -132 -1739
rect -65 -1792 -62 -1738
rect 189 -1776 244 -1773
rect -175 -1796 -62 -1792
rect 254 -1791 257 -1727
rect 364 -1732 367 -1662
rect 408 -1711 412 -1506
rect 440 -1512 450 -1507
rect 447 -1600 450 -1512
rect 507 -1521 510 -1430
rect 550 -1445 562 -1440
rect 559 -1466 562 -1445
rect 550 -1471 562 -1466
rect 559 -1541 562 -1471
rect 549 -1546 562 -1541
rect 469 -1551 492 -1547
rect 559 -1600 562 -1546
rect 447 -1603 596 -1600
rect 541 -1612 565 -1609
rect 541 -1615 544 -1612
rect 442 -1618 544 -1615
rect 442 -1622 446 -1618
rect 408 -1714 438 -1711
rect 434 -1718 438 -1714
rect 483 -1723 486 -1698
rect 541 -1712 544 -1618
rect 593 -1631 596 -1603
rect 584 -1636 596 -1631
rect 593 -1657 596 -1636
rect 584 -1662 596 -1657
rect 471 -1727 486 -1723
rect 354 -1737 367 -1732
rect 274 -1742 297 -1738
rect 364 -1791 367 -1737
rect 418 -1776 473 -1773
rect 254 -1795 367 -1791
rect 483 -1791 486 -1727
rect 593 -1732 596 -1662
rect 647 -1708 651 -1503
rect 679 -1509 689 -1504
rect 686 -1597 689 -1509
rect 746 -1518 749 -1427
rect 789 -1442 801 -1437
rect 798 -1463 801 -1442
rect 789 -1468 801 -1463
rect 798 -1538 801 -1468
rect 788 -1543 801 -1538
rect 708 -1548 731 -1544
rect 798 -1597 801 -1543
rect 686 -1600 835 -1597
rect 780 -1609 804 -1606
rect 780 -1612 783 -1609
rect 681 -1615 783 -1612
rect 681 -1619 685 -1615
rect 647 -1711 677 -1708
rect 673 -1715 677 -1711
rect 722 -1720 725 -1695
rect 780 -1709 783 -1615
rect 832 -1628 835 -1600
rect 823 -1633 835 -1628
rect 832 -1654 835 -1633
rect 823 -1659 835 -1654
rect 710 -1724 725 -1720
rect 583 -1737 596 -1732
rect 503 -1742 526 -1738
rect 593 -1791 596 -1737
rect 657 -1773 712 -1770
rect 483 -1795 596 -1791
rect 722 -1788 725 -1724
rect 832 -1729 835 -1659
rect 822 -1734 835 -1729
rect 742 -1739 765 -1735
rect 832 -1788 835 -1734
rect 722 -1792 835 -1788
rect -65 -1802 -62 -1796
rect 364 -1801 367 -1795
rect 593 -1798 596 -1795
rect 832 -1798 835 -1792
rect 593 -1801 994 -1798
rect 168 -1802 596 -1801
rect -258 -1804 596 -1802
rect -258 -1805 171 -1804
rect -309 -1878 -79 -1875
rect -73 -1878 159 -1875
rect 165 -1878 403 -1875
rect 409 -1878 596 -1875
rect 46 -1903 49 -1888
rect 284 -1903 287 -1888
rect 434 -1895 528 -1892
rect -48 -1906 49 -1903
rect -53 -2190 -49 -1985
rect -21 -1991 -11 -1986
rect -14 -2079 -11 -1991
rect 46 -2000 49 -1906
rect 190 -1906 287 -1903
rect 89 -1924 101 -1919
rect 98 -1945 101 -1924
rect 89 -1950 101 -1945
rect 98 -2020 101 -1950
rect 88 -2025 101 -2020
rect 8 -2030 31 -2026
rect 98 -2079 101 -2025
rect -14 -2082 135 -2079
rect 80 -2091 104 -2088
rect 80 -2094 83 -2091
rect -19 -2097 83 -2094
rect -19 -2101 -15 -2097
rect -53 -2193 -23 -2190
rect -27 -2197 -23 -2193
rect 22 -2202 25 -2177
rect 80 -2191 83 -2097
rect 132 -2110 135 -2082
rect 123 -2115 135 -2110
rect 132 -2136 135 -2115
rect 123 -2141 135 -2136
rect 10 -2206 25 -2202
rect -43 -2255 12 -2252
rect 22 -2270 25 -2206
rect 132 -2211 135 -2141
rect 185 -2190 189 -1985
rect 217 -1991 227 -1986
rect 224 -2079 227 -1991
rect 284 -2000 287 -1906
rect 327 -1924 339 -1919
rect 336 -1945 339 -1924
rect 327 -1950 339 -1945
rect 336 -2020 339 -1950
rect 326 -2025 339 -2020
rect 246 -2030 269 -2026
rect 336 -2079 339 -2025
rect 224 -2082 373 -2079
rect 318 -2091 342 -2088
rect 318 -2094 321 -2091
rect 219 -2097 321 -2094
rect 219 -2101 223 -2097
rect 185 -2193 215 -2190
rect 211 -2197 215 -2193
rect 260 -2202 263 -2177
rect 318 -2191 321 -2097
rect 370 -2110 373 -2082
rect 361 -2115 373 -2110
rect 370 -2136 373 -2115
rect 429 -2130 433 -1974
rect 461 -1980 471 -1975
rect 468 -2068 471 -1980
rect 528 -1989 531 -1897
rect 627 -1903 718 -1900
rect 571 -1913 583 -1908
rect 580 -1934 583 -1913
rect 571 -1939 583 -1934
rect 580 -2009 583 -1939
rect 570 -2014 583 -2009
rect 490 -2019 513 -2015
rect 580 -2068 583 -2014
rect 468 -2071 583 -2068
rect 361 -2141 373 -2136
rect 248 -2206 263 -2202
rect 122 -2216 135 -2211
rect 42 -2221 65 -2217
rect 132 -2270 135 -2216
rect 195 -2255 250 -2252
rect 22 -2274 135 -2270
rect 260 -2270 263 -2206
rect 370 -2211 373 -2141
rect 360 -2216 373 -2211
rect 280 -2221 303 -2217
rect 370 -2270 373 -2216
rect 260 -2274 373 -2270
rect 132 -2280 135 -2274
rect 370 -2277 373 -2274
rect 580 -2277 583 -2071
rect 622 -2187 626 -1982
rect 654 -1988 664 -1983
rect 661 -2076 664 -1988
rect 721 -1997 724 -1906
rect 764 -1921 776 -1916
rect 773 -1942 776 -1921
rect 764 -1947 776 -1942
rect 773 -2017 776 -1947
rect 763 -2022 776 -2017
rect 683 -2027 706 -2023
rect 773 -2076 776 -2022
rect 661 -2079 810 -2076
rect 755 -2088 779 -2085
rect 755 -2091 758 -2088
rect 656 -2094 758 -2091
rect 656 -2098 660 -2094
rect 622 -2190 652 -2187
rect 648 -2194 652 -2190
rect 697 -2199 700 -2174
rect 755 -2188 758 -2094
rect 807 -2107 810 -2079
rect 798 -2112 810 -2107
rect 807 -2133 810 -2112
rect 798 -2138 810 -2133
rect 685 -2203 700 -2199
rect 632 -2252 687 -2249
rect 697 -2267 700 -2203
rect 807 -2208 810 -2138
rect 797 -2213 810 -2208
rect 717 -2218 740 -2214
rect 807 -2267 810 -2213
rect 697 -2271 810 -2267
rect 807 -2277 810 -2271
rect 370 -2280 992 -2277
rect 132 -2283 373 -2280
<< m3contact >>
rect 593 -994 602 -989
rect 776 -1001 786 -993
rect -154 -1431 -146 -1425
rect 275 -1430 283 -1424
rect 528 -1897 533 -1892
rect 718 -1906 726 -1900
<< m123contact >>
rect 529 -844 536 -837
rect 550 -842 557 -835
rect 750 -855 760 -847
rect 522 -1371 535 -1361
rect -159 -1414 -146 -1408
rect 270 -1413 283 -1407
rect 499 -1413 512 -1407
rect 738 -1412 745 -1406
rect 516 -1421 522 -1416
rect 562 -1422 572 -1417
rect 755 -1418 765 -1410
rect 800 -1419 812 -1414
rect 504 -1430 512 -1424
rect 743 -1427 751 -1421
rect 677 -1810 682 -1805
rect 586 -1820 591 -1815
rect 526 -1871 531 -1866
rect 713 -1891 720 -1885
rect 730 -1897 736 -1892
rect 776 -1898 786 -1893
<< metal3 >>
rect 529 -1361 533 -844
rect 550 -1406 553 -842
rect 518 -1409 553 -1406
rect 596 -1409 600 -994
rect 753 -998 757 -855
rect 753 -1002 761 -998
rect -152 -1425 -148 -1414
rect 277 -1424 281 -1413
rect 506 -1424 510 -1413
rect 518 -1416 522 -1409
rect 565 -1412 600 -1409
rect 565 -1417 569 -1412
rect 745 -1421 749 -1406
rect 757 -1410 761 -1002
rect 779 -1406 783 -1001
rect 779 -1409 808 -1406
rect 804 -1414 808 -1409
rect 682 -1808 758 -1805
rect 591 -1818 736 -1815
rect 528 -1892 531 -1871
rect 720 -1900 724 -1885
rect 732 -1892 736 -1818
rect 754 -1885 758 -1808
rect 754 -1888 783 -1885
rect 779 -1893 783 -1888
<< labels >>
rlabel metal1 11 -680 12 -679 1 A3
rlabel metal1 11 -688 12 -687 1 A2
rlabel metal1 11 -696 12 -695 1 A1
rlabel metal1 11 -704 12 -703 1 A0
rlabel metal1 11 -714 12 -713 1 B3
rlabel metal1 11 -722 12 -721 1 B2
rlabel metal1 11 -730 12 -729 1 B1
rlabel metal1 11 -738 12 -737 1 B0
flabel space 56 -748 57 -747 1 FreeSans 44 0 0 0 and1
flabel space 118 -748 119 -747 1 FreeSans 44 0 0 0 and2
flabel space 178 -748 179 -747 1 FreeSans 44 0 0 0 and3
flabel space 238 -748 239 -747 1 FreeSans 44 0 0 0 and4
flabel space 298 -748 299 -747 1 FreeSans 44 0 0 0 and5
flabel space 358 -748 359 -747 1 FreeSans 44 0 0 0 and6
flabel space 418 -748 419 -747 1 FreeSans 44 0 0 0 and7
flabel space 478 -748 479 -747 1 FreeSans 44 0 0 0 and8
flabel space 538 -748 539 -747 1 FreeSans 44 0 0 0 and9
flabel space 598 -748 599 -747 1 FreeSans 44 0 0 0 and10
flabel space 658 -748 659 -747 1 FreeSans 44 0 0 0 and11
flabel space 718 -748 719 -747 1 FreeSans 44 0 0 0 and12
flabel space 778 -748 779 -747 1 FreeSans 44 0 0 0 and13
flabel space 838 -748 839 -747 1 FreeSans 44 0 0 0 and14
flabel space 898 -748 899 -747 1 FreeSans 44 0 0 0 and15
flabel space 958 -748 959 -747 1 FreeSans 44 0 0 0 and16
flabel space 850 -852 851 -851 1 FreeSans 44 0 0 0 HA4
flabel space 667 -852 668 -851 1 FreeSans 44 0 0 0 HA3
flabel metal2 780 -990 782 -989 1 FreeSans 44 0 0 0 L7
flabel space 430 -848 431 -847 1 FreeSans 44 0 0 0 HA2
flabel metal2 598 -989 600 -988 1 FreeSans 44 0 0 0 L5
flabel metal2 361 -985 363 -984 1 FreeSans 44 0 0 0 L3
flabel metal1 741 -1043 743 -1042 1 FreeSans 44 0 0 0 L6
flabel metal1 504 -1039 506 -1038 1 FreeSans 44 0 0 0 L4
flabel metal1 39 -835 41 -834 1 FreeSans 44 0 0 0 O1
flabel metal1 98 -835 100 -834 1 FreeSans 44 0 0 0 O2
flabel metal1 159 -835 161 -834 1 FreeSans 44 0 0 0 O3
flabel metal1 218 -835 220 -834 1 FreeSans 44 0 0 0 O4
flabel metal1 278 -835 280 -834 1 FreeSans 44 0 0 0 O5
flabel metal1 338 -835 340 -834 1 FreeSans 44 0 0 0 O6
flabel metal1 398 -834 400 -833 1 FreeSans 44 0 0 0 O7
flabel metal1 459 -835 461 -834 1 FreeSans 44 0 0 0 O8
flabel metal1 518 -835 520 -834 1 FreeSans 44 0 0 0 O9
flabel metal1 578 -835 580 -834 1 FreeSans 44 0 0 0 O10
flabel metal1 638 -834 640 -833 1 FreeSans 44 0 0 0 O11
flabel metal1 699 -834 701 -833 1 FreeSans 44 0 0 0 O12
flabel metal1 758 -835 760 -834 1 FreeSans 44 0 0 0 O13
flabel metal1 818 -834 820 -833 1 FreeSans 44 0 0 0 O14
flabel metal1 878 -835 880 -834 1 FreeSans 44 0 0 0 O15
flabel metal1 997 -750 999 -748 7 FreeSans 44 0 0 0 VDD
flabel space 142 -874 144 -872 1 FreeSans 44 0 0 0 FA1
flabel metal1 45 -1246 46 -1244 1 FreeSans 44 0 0 0 L1
flabel metal2 -309 -833 -306 -827 3 FreeSans 89 0 0 0 GND
flabel metal1 193 -1250 194 -1249 1 FreeSans 44 0 0 0 L2
flabel metal1 923 -2355 924 -2353 1 FreeSans 89 0 0 0 P1
flabel metal1 939 -2356 941 -2354 1 FreeSans 89 0 0 0 P0
flabel metal1 825 -2354 826 -2353 1 FreeSans 89 0 0 0 P2
flabel metal1 573 -2355 575 -2354 1 FreeSans 89 0 0 0 P4
flabel metal1 801 -2357 803 -2356 1 FreeSans 89 0 0 0 P3
flabel metal1 126 -2359 127 -2358 1 FreeSans 89 0 0 0 P5
flabel space 75 -1902 77 -1899 1 FreeSans 89 0 0 0 FA9
flabel metal1 -217 -2340 -217 -2339 1 FreeSans 89 0 0 0 C5
flabel metal1 -120 -2339 -119 -2338 1 FreeSans 89 0 0 0 P6
flabel metal1 -22 -2274 -21 -2273 1 FreeSans 44 0 0 0 M7
flabel metal1 216 -2274 217 -2273 1 FreeSans 44 0 0 0 M8
flabel metal1 364 -2289 365 -2288 1 FreeSans 44 0 0 0 M9
flabel space 313 -1902 315 -1899 1 FreeSans 44 0 0 0 FA10
flabel metal1 439 -1795 440 -1794 1 FreeSans 44 0 0 0 M3
flabel space 536 -1423 538 -1421 1 FreeSans 44 0 0 0 FA7
flabel space 574 -1890 575 -1889 1 FreeSans 44 0 0 0 HA11
flabel metal2 429 -2015 430 -2014 1 FreeSans 44 0 0 0 M10
flabel metal1 653 -2271 654 -2270 1 FreeSans 44 0 0 0 M11
flabel metal1 587 -1810 588 -1809 1 FreeSans 44 0 0 0 M4
flabel space 750 -1899 752 -1897 1 FreeSans 44 0 0 0 FA12
flabel space -122 -1424 -120 -1422 1 FreeSans 44 0 0 0 FA5
flabel metal1 210 -1795 211 -1793 1 FreeSans 44 0 0 0 M1
flabel metal1 358 -1817 359 -1815 1 FreeSans 44 0 0 0 M2
flabel space 307 -1423 309 -1421 1 FreeSans 44 0 0 0 FA6
flabel metal1 678 -1792 679 -1791 1 FreeSans 44 0 0 0 M5
flabel space 775 -1420 777 -1418 1 FreeSans 44 0 0 0 FA8
<< end >>
